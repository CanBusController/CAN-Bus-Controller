// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:39:00 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
M7Zl0KOG+hpgNcQCL7hf+fWcQ311/1kUJbPyBXKtNbquNyMYxN1fNh5i1Lx4m7DN
LdiznIaw3xiSCwG2TlNpPyJHaiijgz08tmy42FJyJzgRNidTHiOGgkjiNcBQRQ1A
f2DpzBy3ZBwmLeJLI8EM7Blk3KFW/f4hi8fekD2G7mg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11808)
EJKQ57jhocZ/1E+QbNEkt7bP8lZyqqi8w2NK0HUXcWSAO7hcqsxo/BC2SChAzpAb
GRY+djqp86kFr0ovHp6lIWoYZBp58QuhIbIka2VNHtbq5ig6iMsOWME1Npcxw0C+
PvIK+yPYB/ULDLmTWbG9YfSFdlg109PC6ajJYVVx2igLQdI+ChaN3rRODZWHmwnB
b8sJPGnrFYZouYl0NZJUbi8NFxkuTHbRGPWiAGQJrRopE+lItfRFS+mLeqW2iLvN
cpiLvpWA5h/3+oVpe4/kmh/QoAX5rVW6CAHePHo1/VwyLpnmcrNaFNbICOJxvlhJ
XgQ1VsduUCPNRtmqFU6KUOFUhT53j6nCwqSsoZM6/895WzfhGJY017Nqb6nQ91da
LeBFaVBW4LG+S6m2h8AXkEvgicEZ7FDZ/gPx2Zj4Sa8kVUY4+gd0f4qEY5GMTeAf
bL0WBlssd8FPoWnSt/yQEpgfJ+QAc7j53Fwoc22uaRscWPfAf7UBm9ZE2IEVwipP
ypXkENLvjAoH3r1ysCWq3bwEH+zWoV1HyVsp/dw6hJX92XdPZ/5jnoeHlKwLRaqd
hJKHgqH9syTYHbtU5I2JEJJQjnLIqP+6jf/DbniE13ql2KZn8oaqC6VknPj8iC+m
OHfX0h4lkaF6kwwOtify8H+bo8QTOBxw4UCo2Hkh3f10wacqWVgBZNwH/3h1Q8lY
TBEJCep1gpTKMKURmOnA5Hvb8MghRwGfftwoXXe+4THiYsSEOCc9OrFTkcsDotxF
vwQYQGgzGYHtl7ZGeAhB0DNIjytEYojYdZdADnF2hjgSytoGXlEVXSpebHuR5l1f
xXQmWC/B1Z430Eg6L7NEfoqDa1jr10716g5kRhU4/ddhBpgJ08Dt2Wa6Hl7rXyLL
17jdRGMFEl03rT6WbQkrO5F6YxyYndwTbYNAomD0Px4QO+8xye4F1McbS9OR96T0
+nWzFSLWf63IKCSY564eHp1KPX0yT0FqFXTgrqi/shXlMyiqAJfXaRHV3CZkeHXu
IXeM2ZRVV2PoDvbIOoShd5BqRGziUZwB2H4T2jtcZQ8punzlegJp8+clCq1lw8s7
/EKFTQAZp9ZlZsUsfZVDGIoRZMWXn9l3aNCqEAI7WFvvs8oq94Eccn46cvkyzt5A
/PoV4j1+/abfUTShYT5yNmLkPy+FYC2SjC7ifNgVHF4x5UoCXFsdJbbpQH/QhMB+
kfPDvMjn3zRsmfG65s3Pus40xBF+n5UhZepwwg8xHrEUbtM1pPjo6d5Tdy+hlS7t
zW8mPEiPaYlltcvdbw50YICC/ZKDFsA1sm1W9hRGaqBYgNOI+5tSCl13scnYCX2c
E8qSVAluaq98QOrJVd/BKYonKNxMyzUsvDFy7JjwwL4SKrq4ldGedGt6qj45HGi6
XpczzhWUzgXqQ/aiBBv/fqIv0tDqg1WQ73puFCvyik5bla3x8QOTKifwz5eUCrdq
hRD3D0BpA+rR0/N+Q8EIGga4Xb8jZLYCYNoG7m5VN65PhlNmLRbjnVbwooyT2UzQ
NGU6Pd/0g6NwqH4+qSgYHoawqiZSC6R3QauZNO0/F6rxE+XaaoSwVOPi+7gZMjx0
kmqRRJXb9ED67D2aA2+0Tly1IDH6pC/FI/+H2ve1JQjWMnsFE4LkGdcvHO6bTb+u
zGsC8/sqXoFDy2C2WUf6aXs6wzt/fKbh44OJd1N4nt7iccI0u3hKvABEe3CHuNwE
8A5KZM5k5j3BgJ9T6cSHqfe03DaDgsqMSTZ2lUGkgc8fWujLnerxMHBfYHX+Ptav
bN/QE+8+z/F9aSCqq7Q1hJl+eELhjQmeei/qiFMR22MR5egVwoYN0xGTXv7xDuk6
18EsrO7XIa8ALge5fsAGJoYtshu08fI750nEssIRFNe/sLU0OytOOujPDd4g7vXK
rqfZicO9d/xyy60bee9F5wACsu+g2nI5O86DVN3n0fVkpQtPVqLzxwsK+Mvk6Oab
l7swT9xq7OnYlaLnGt3gGHb+c9shrAblWES+xDoco0S55OASnXfw8B/GIuqSBuy/
ljV7dtZAA0k7F9UmCa56jklx+7Z5qsClTQXfz/nAYobYCr9E2KZsN4gOMdIxyLJc
KnCmPzoLL2tSlSueTs+zljdX7L3zZoSR+OjBAgxTBqhggPksB/ap5FxDjmWHLEjZ
7ur/K+NINdWdL0WVRHRDN9pwsHr6HpKTSPZSMJZGzKT2CUrEQyOSHyC93K6kC3ev
/Kpbch/DlpXMT+dh0cDXAuvTeBuIym4gYtMdD9YtsCSPaEMI/ahXDGHQAjHKnEZL
benSSYvCc1p56kjNiK1RB8FmMm/F6Q+Ft3+gv80uApcWrLbe6sLAjRRgNe4tioiZ
ibANyeacgEm/us7SQiNHCZO18SDkXLzPJ7FSBPYaZINDwONhRuYlMqtV7V2n1Ik5
MgCAXCksBb7t+8gN9jgAWGDE1dM3nJQ0azn6f+ytdjYkd1cBdm3gBgZ/42eSP10t
//VoyCjO0NKW1ThHB/TKY2NhYamnl6n7xwyUEiyajn1TpLCFY+L+BJrBswF+o0WK
rRUQJbAr1HthPJTgOF0/OboR7RBitX8uYFt2/A8EgWDnLPtS4cRFwOnAUOTwAwjG
0xxdy2x3qRwIXjHn9rfXiCC8PmqJBYJEH1vqBwmfdM8xfNwuIX3h5v1zxUFfSUZG
UEWGP59lDs959p1HIzYWTpqdHHhQ2XeRWcviXPPVrNsVZzN6p+/DDOL8l2ZrO+Qs
KclxdV9J2nEzm7f+FqbVzcenRrGowvl46V/bC9hHerW0bmjwtfxXdkHRrAgqu0GY
4Kf8sJZdqCgYB0JVeMvZsod0Ts3Y4jInhYAkantmcK7bd3a96mggSu3X5GXd+juX
6f9QwvEtkTrfIPvIqXjYo+QIoCpRCgoe6LlLTAFiPoAeofzhkSl2p+8dNmwzkAGQ
QXv3Z5tGkRVFlp+kpV/ttSlo2pzXcE2jfuSqz3fMuK2uQw1ydB5XS13tnROfBtkB
BBawGW+m6cH9gwWBVReeyCUKYc67dz6oh6V5XCO3SX9B4SEwKELej5U5KOn5y2Vt
Ts3/6ljDdsF436baw2vjVaU5ZSNPshBpRR83cDxwyGtWHRhyfCTzAE1Adp4Cx+tq
ijECZoHr2+eEZhxw0MnOhaDOSGx5Yxu+aN3VMHoIrCRL7cExpkjtNX7DXfYPljDu
mWfZazTB3K7JQXIrkGCLFAmexMDXR4bEfLTn1+l7DpTsgx30boee6GKEwt7DRj96
P5WcLBoAaUpNIDWKhwKYQvYIAGgMAC42mMFlN6JGlLIuROa33rbwuXt3Cm5TuTPC
afKRBDZYt04nk9JG2TuGyu/mdDLGBanQbg56/Y/PIZ4F/HwlVh8IPqOg+yef0tbi
/iBUx5xAUM9Rr23dX09g4NMmm7WLCczb1U4R4SV9yuk4Fq/I1HrXkjJQEde1TbEK
mVa4ppKGnwGI8F/oZ5gEjlK6Or1sOafTj41DZv+khpM6ob98lUsFftIEIo0ejmkU
5XFGSqdECgjs7XO9Azy80k2s8loS/CKoAU+Yybidk8U44Kcz62cbPKobeR2Ay9wk
kaL+0N5SW+BPINKbggNEy3IRh0B9ElIJ6FCIPCEC744eFs882LL7eAsDLpIvYFkh
YkXnUzN6k1jxniVcoOJjWs5k62oQgm64T4W8raCaqOpQ3MLqbnNUXufZfX5TJhzm
MUm+xnlqCyMvo5MLV6LXEn5JxC3QYinM6nA7W0SbZVLFvOYyVPSaD8JZ7LBWoqKB
WOM7YYl2VlbfLhCpLcl86O0Ce6TLl4AoHBcROyRO1RaFK6QX3cpuzl9jCgMoPf0s
46R/k3/CR4sudC1GxWQMougXN+p4R6FaflEdi38siPRFFzsF4vrrY4P9ywgsN6Md
L21PWwnyB9a9U7A7sASHpr6lyBO7ogkorBcPT3uv7bGskfNGzVWQ8pmz2OPKWWVg
4aeF8XX7wakWR3iFPGJvHrFiNg8JzSB5lxTk2WLpPm+rKSOFSMF5yR6T0rnOeFz8
/QKV2JaEan5BTiVaJUETI4ddQAA4v6gbCN18kicMfhT9swtg5bSkmc/dRLMLufP+
RCwB+ucLdj//i8NIG5VrDUkwJ3Ah59FJ/aZeB/yDnj6U153Eb6xF804WbeLrzdLX
iEf0VZ+Y+DlQ0gktIBtWkTuBRY7PTZmTWMrbyrjiv9wihNaZrXgXyDQuSRlkt9fX
r4Po+Xq3uYyJyl0rb8nI9YvPGolqAngsSzRTNlX6NNntBot0KZ8l3WWbNcUyywLF
8c/rzglSqnB0kTOvfOidtRGo4wSzZup1vNNEAYI/zTQW0Ux7RCTyGdl5LcOwdr6F
T9V2i9ik7G9OPp9QCtDzrtYlyBVy6vQqV5UQEwjswmCfXv6rtN6RWU1nH1o69W+U
JjGqgVIq16kVoKAHmT9QM0fkIlz0Wa6ydwdxhqQC/g7bWNUDmh9gOoZlIamlWruO
qRlgn8gzNngQq7c+HrcnmnCJXKFEouoxWNGj6jYcKTrGBHCwFrJIMwFsavUjms3T
Ag3aClSjD7zQ292FOwwVe0I/MhbJ3DHrMF52jBeLfObX5CFgILj0RkeNWCHrwFh8
JhS6bpVPmd4u6JExSgviFh9ayJEJXE1sNVxLuxYSEJPkPI4K9u8d8EVjyTQ1TE39
YLdj+kBZLogCx9QGGS15cW9qCC+T0gC4TFGoHhiFxi1KalV6t+ZyXllKJNar1nef
kwqmxmJ4NWOJRI1/PeX2Z47nuFgW8sLx7qzkIB9V05NpzM/G9uBrfKtCQWbSjqqH
zA/2UMevFVKtFRpqU7TLuces1CsAMPa/7qAYyBu2I9xjxjSLs9tm3MrB1+CNkXC2
SIPxE2i0IVTl+Eahk47WDaPmvaljSDKHC1HNPvaxJu6kjZgL2FcmVHfS4yI/Su4J
Lo2xiAnpkq2nyCLCNeMru1cI/vyl9wgJ6Vo4IUxisGo2zbg3rql91mbpusz58cVK
ZGZc3Evih953xZiiz2XjduX5QYW8JtmmFn7GiVkP5g9SXefTvioNDzp0hj3Auu7+
AlqOiJqc+F1DeM6bKh+3T7VFbKe6K9u0Axj0mkfiIa2/X2qmk/20sbNXjmxd7zVI
Sa1n5w0QQNtB5QVh2zjP/UEZV0Q+JDl176GzwZPg11jy6WuJty28npzUXTgXiNfo
rgF4hbB01Aq3/CzEJTnYcN1rCV8vx8vU1VHHw7cMaFB+Xu0+mPyALxUywy28Ua/o
iqygLv0D92KZHTv4KJbjVeWdu98BVRMJHMJUjGl0nrYSKaVVcXAAdto+1JFniYZI
ZB8132C+rFGQSU4lOkj06ytaQad/N6tx3m7IJHT/A8K9Y0wZuwanhUhQCQvO6aol
mj/higR8ecOzQLDVeWxum1YnpTEAcl6xHLMyRfDZaJDDlQxVdK8oZGTv0/qLcxb9
DLI9RSWy1LRj9nOofdecrgLK8B8ohk5MfaWaZw+1FCRXSnq+25cfVcMhQaj3tDfm
hDemPFxZE8aEQ49yipzu51vyFdNiHhbkFxsFGfSFIHriBatPjRFpnbOFkoO5/t5V
4ywBnKPrLWTj1RrTOBoCTcWpcfED4uNQQUAFoAeZ+gBygm7b664P3cDjUQpDAYzh
/nOxovy5UFpPWzQYKpLvpP9MiVPjrQE4XxiF+X9h8lfKvzTLVmmbzTJ+KyZtsf5m
bBhNekcfR+6YFCmAV5aDtUbPZGVE4F2OPY524NXJjVxJCIo6Cm4HYjYFimRNOU1s
HNN58O9ela6DbK4rJ63EyjWZVOqbN4IKkh9J7sfJmUvlSe/GkbjRZtHT51HBxVzK
yNdWFTHRADWjXthqothWb1gyBWS4nMK10sI4g+1xsaHwCTfS+gNnj3NX6QxtF+hP
Ca+SnUJfqYAINt31Wowp7QSoxi4FLLXSWAqhVkUM2hvNbHgpCGBeNAYSFjZTYm5A
ffMUceGbg/PU38FGqUj3vgqTdSmsYjJ//tXCRIuy8KlP0Wi3OGSSkh6NildjLCVn
nTw0d3O5XmiAuVsIYrBFP2PFASWqgYnAtiHGD2F4DOBT3YhNyzBZzqRyQqPM4dIs
QrO5zgiK3/ddCCjGjbpfjJeSC5wsB7xGlYAhJQ9VCbEBUos6TVvZfpuZB42IKzPG
tuaYWv/t0gOOL9/4rZCUi4GKZ7NC33RUdJLtuV028DpR9sNDH0NdkutpgSePcUxN
In3v4ggSpc2YeXqi89sxSWl49Kcs/Cu2ClnjRmKCTWrtE7Rr2mM85aSuK0HVHId/
VzGev0i4AZXIAYlHNSp4X88Eh7c5LZub4IHllXswY09Q5q5W6tzog8VfQCQ6a6yY
8r/dBJhOl+JLpG73humagjz0aFQFL8o7CK6Ke2zmgJKQxCpaxcLnCwRlIXZK1jqO
P9HBKgIHXGMSRnlvFOPDyRQGXUubyaABrbadWJetytW4nUH6wmcBQWNxpzsBq+Ns
X1F0dKXz1xSx+yBtdfCETxlUO1f0+S7FCn3VNfsy0qwaKSNsDraz7L33wVbT+Y8Y
BZgqRGzP3WgFc/B2TRFqp3l2rOyx5L1LzzU20mBPGithXSObDCaFiM6T9ZZ1WCFN
NPXmEWhBbJaYTwrsy5h4LQQedLQ53/40upJzH6zce3CGcFSLCf7Xqh9spBHyz6tF
8I6qMPnFvpNu26G5LxMKJp0T2e8d/malnfdq1lAUIG2UypBWae0FYtT/0B6xXJAY
aumHR7BgJlvwte+KSj/zb7WRfjn4Pdy0GxycG1W4FpN+S8fhu71WuWiOFJYQ0fXG
bwZ1Z/1kuzfJsluQDJ2gpULh1xeJg3Nkm/8nwAkXKW2hVLtczzneJR3wx4aBLYsj
pA3RdzK+dhqWtxKxWXjkI2+eX0xKujR4n7nnkD+3J13G5oVCrX8vz1u7ADoxIJXa
JzCc4ao0GQ7N6+kZ2umvUmrY/vf7LDrwdwsCJDiauoZI3rfKT5Va4hpcCijaaRqH
eSuVv95DhsiIEGfEFKkXyzlkLjeiIWEvZyg6+YoZTCmQF92zEia3N29uJYwt6sii
FCFkB/RiqueuchdEevZuxkpaw+zPAMGUFgyOrUJ2NnxQArpwekQzHm/rPK3ec9T4
MbCqu+fKEvexXFilGPjyAh2pCGE/kME0y9MdQfnUKJTyrCFKAMtA2dtXxKMFhDjR
GpMkyBV7k96CFs4Diw0ntk6JqzTS6BgKCVQpt4p1PqFYbT6J+/QgJmWzhnYQLpEW
PLFeV0uZzlEPe7m1JVg4poPLEKD5hFt+8w5iWt1L/ZfcPioAX/Ld/CkRnIp0eKjl
0uT98Hv+IGPSfVdU2iZ+pT6REvXxg2+blzQIAVh5VsVv3LRVCzTAgWjRHIRt1HKu
9IQKgiyRYCB4GLGwV+M2ftXf8aTicxA1aRoNMdGMct+9rYEitTnZOnm1zMJLXyH7
Ms6X6wUci3vIW55KSvQQeZ/+LcYRIO7oGmYdncMVOxaUrASIYVfHbAI681UKZa73
6Qzxpo1lcZwxbK2qJhVuqoZnIVhr8fMT3ut98mh4xE1icsA18vuyMLJCDS4i8FY7
+fIBfgSSSZh2L6BuN8+BckJvMGm57eIl2a5Y7stpB2eVpqcl21clUKeal5ZTSJg2
OfqlBWfPHtzgu3ir+91eCn63xjTzySIchGVaKcELIrg/O6zUexUxJtoUqakSEKA4
zYbJzWJ/Xwxh450nm2e/SrcG23lh7Gyin/i+VbfR6cfxXkiWsYuFnCbcIFKrQn6r
nLQy+z6uz8pqPPZ/PMFTTrBJLbHE/AAMsEq3f6NV84V94UYGc/kU39cgEABjbcC6
NrXkTM1RNLgTmO5fZ3TtQH08z/az8+Ir4V/dH9IzZUCx66+69LOAQUc65JiFLkvu
xOVgsHHl6CctIcaS2v/NQM8nC43HN3PFl4xudzHquGFN2k9Ff90WOSYHc48CHhxf
4SmQwbwDYLwCzQI9JGCTzK3Zmaju9udU6SnFPbrnsW1DbDbFVeFoXT4BQQSVFYln
xfKKC+Kd7yk/sN44P7KCglKIZtVTqNES1VpWwU5eu2F1eXZ2+JkWO2v9fJ6T2pgu
KMa8KSRj/OqGTGa1ZVD4FYDQqJDbzZ78GTIB+JNhhFeVIJWTEhQ9K7EHPVAsC9K0
yu2HoKmKwAQYEoW2rFsmaLCtAvdJeSLXWRmfA2lBJoM/MH12SL9Ccu8jgIxfsxYS
7cus3ww20bPGBV/5FXdY5nlDgI5QZ7BeaasvOdqDmwDPcgOz+3+R9dd8pifHTFWv
ckozYkNKQOozPRw9dMmTgMt33YWJl+sOUILxM3muIKbzrvJcs14jQfreao9dX/W8
Qwt1vcakLNDOXmr+I5oQcOghb5PZvLtZif5auBrH4MCD1O41rUHDmDkBWczsFtqc
xnvy5CqBOdOu9mjcJ8MnB+PhWuVmLW+GACES8Ou2+q+L2pJ6sb04JlBWeqFD6VCO
dgRmQ1+rT21XQj8nnIY/oXDh1KTcSgQBz2W1onmgnCOQSrc1m7tiH6B8g4rgQ5Ag
ybUWdOhL3gdJhOOT1cbhWqCEO/dWa9TkdagCNd1t4FgWFOYCj3qeAUPNSWKeYyt1
q2hzINzW0MD47K0JIp3SZOsExHNB35fjWFTHDEkh+PqkGkTvq4TZciVA/WAB92L1
2IJTSz53VKrl9TbSo+E9zlMFnjZ63fBbhrzaIVk14aB6S1TMbRQs7DOJ3i529TWX
OW28s7N22/6mFqaVRa5hnhAtkjr6XVjKhh6vrAQExXOcPgcU+p+Dru4eFz5lj8QJ
HwY4KcW9bGAf2mvw5sym7LSfDV6gElLCQtJrNPbdT15UEusR0BMhOXOd95FrZDkh
XW32+S4T2S72dSX86VNQcq5ygRITbXeRGxEls5bnifgnWZdqC/8bL5cs9i+AUcqH
lXLsStFtSa1+e2rVfjNU4gWiXhPEUu2tlCWErxRdVZJ4qyu1qZqkYh0gJus92QFr
VjkX3jLnQjwqf+tBA9LmvL1MCsYAmqTlgLmSvyw4vwFuHi/uBqPkG8UaHuzoqGli
PUJz/+7uYYr7UgpX+5MRzROXmmfJPdrM3SUS8SuGoYVq/4i0AtbdCEUvkIxB561Q
wh8JG//wUManXboMl2JW8O2ZLORI9qIYSz9dYVNGs/RH3dJFulOHsxesDVJm0Lzg
p6C6xgt9H48o1+8UVMD9GGVPMK4l+kfy+RcsKldyOzrLhCV2iZ4/VDBjipLRxSnT
KVff/Z1KB/jg+Ui9b5mPaKe/hzSf8JSzzOM2na9mjsrHv1aGMwc4rjRXAcyQmj9N
IXcbH6kCSA33UQt5+f+NrKAdqQoIQX3tiLd5DUVTKuECSn2CrMD+uheShpcvLMxR
nYerRzTlDAivcpFU6OcI6utgRrjEoeZ63d8a/GJO2VPFg84gz6Y5Tsc0Fmxpr581
ufOfkToldK5l9B3jvlg/RUK0NOj5vqo6YzMN5fAB1GxA0TU5ET++q2ZqVRBDgK7D
GuyhRKYhYJgwg+5G37xRBtSyeRmraRp+VHZ+lZJkvhLF2hSggw/bYK6v4a8HYo3f
ZyxOrS7wOFwwE0x1mGGLJ900/ftbyLFyBF75UXTH6GXlxLYckS9HDwTpsUVHXf/n
Td6AUvW9ng9EDGqIvlPM8rYgqv7ag/6QllzKa2gcwleVY6TrhBXz0SL8XV968QdG
K3bI0A8NRJLLtJdWkWdTCkN9A8+oFnX1mhJMC9mHboQSWW9BTErJ3pHkD7wFy50Q
F2Zpe4GXiidMjxuq38FB+ozwc7yktNuQk9XJtCVxvnD5atpMz8AUsoACz931M2vq
jUbJVFr+j98lHOyTWBua/ithZhd4JSV/EBg7ET/7ngijGePrWVc4w83IvYXkjipX
+cdnUZ5TEg62EJ/vgrKodpliRKdCBs66fi9Gyw89Us3+YPKmd+Q4LcDEq9fqdPye
6gESpD2pog2BKyaqwR11Nal7X1fdTkf3druVrcPoQQGoMAUsgrQgdDkKtKMe5L+j
u41E3M+tDrcuz7yfgCYMiwkDaqaTXIrbhgAiZCvR4W4FlIikn0GxmCMseDzScQCQ
KQlWu3nPDvT2o8u9m0VjXMeqS0s96w8Z/rJdCsbgINZk1bu5aqTO5Ax2cCJsz3/l
FZX6PqmzciR4y6X1VkxXDbBBztqM558AFPnqUuwmPQsEaexbrESOBQTmvvTYNize
gk9OZp/hIDoerfGSS/ziNUsNDOn9BMqvf5h3w6imrJcRU4/0L7r9ErT/x7/CF6rR
2H9dq014bSeGq5EMZuqC6s2qsaZA/iyh+GIsFv3ImWRacFArjy6AVIjqNEbtOu98
oFuPlEbXLBz9OtYHmUCwr3z4tmApCUzzD52iXB/5mSBrgRPsWY2zmUDoAJxc/j9V
/swy6s42CMFVj81UWTkZi4m3b8wDeuibjE+CUtXDdVP2wuCilSWV50Dm51gJ9e2c
mFIFIUhOIBFadHGK2VT9muy4QOYjaMGfyZ7d/KbftWgfQXUk/AXACOH2Gj/fkKeF
wBTOYRWdQqEtOTXsLijesN984XUFtW69EZc6rJDh+3ylrGzXqED/AU2mkuiPaeyA
SBO/zTTB6R1P7SZkOPRR9HNaZa2XXqAqL+IsH6P8BthtvgRZJ8xsmcvP8jL3r3ic
+etJsnxV8hnBeVPE1tSObePumyNe+paem/Q6MAmu7Eoe56Xa+947InqMJI2jBkGI
TIeqxWo83XbEgEqdnZxq9C8wxmY402L1gylpwZliyufgduqOLUQ+axiAPa4w6oox
LZTsCrzZjSvKVrbl61qJj6D+Ir1VW06figVclhLf9It4ekqq3fV0tcMPX2mXWGAg
mJKdH3i3T9N8AkPCq0EwqJsYvrRc6PTPDYXZXXUoSPbao52sMbnaa2LPiGJU4jXu
JTX3OULdGpOlhkQZrgpOTUk0r3dru7nrvkB8iFE96FyMEo4KKThJcezDG7TO6eDx
VnjVQU1IZ3k1Skxl+oAgm9WbsIVQKuH8Uxnkgy0maOmZ1xK5TSzRnnZxnvGtQmA+
ffkEMZS2xxd42ZtgYNfV5OjsywIhF49khmdtWLi5MaglcK88lF9eMTbDv4tzaCiX
6cvmVDSoR/WG2v/3vNzPqTedOl+8K79PtrAzNNkhpqI1RIB5hHaaK7BCnN9KVW32
fDx4H1IIPUOLPYMt+DOrQVdOqigX6KOKpeuk4ddeFIVuXPvekr5iEDJtj6gzfXUP
Hym2qBGZbYgLClcaHX3FWHY2bKQs7JRo+hCN0l6zeoY/EwVh/m/DxQq7bmn8Pd70
TLDNiwHgWWioKGawzdgK5GkcoepgMSWcEHdOg2Owfr3PEng/W7C164Nn1uv9ReWk
eIH/j7o3uTdfUNrfu8gajdeBCQ9gxrxIjfkYqE2B4c9GtVja9I5ZEtnphRyd8eIz
XVG+bJTsG82LXeDizoXsddMG+RotK3FxSLiPGbUUPG+ZATqF0p/GdnO8onQgU7E8
5iwiorsttO5VbmBiafAcyKzmxSM4U//09zpgZ8ojW4eIjuKVpa5rcDWjvzP5sVVE
UcXcr3seV6hsd4iPbX260gMYpLcWK/ZEq+r8XgAEIGBXniXhwwlcMyXlwBCDP52g
gnXoVmjhus+/MyqFCk72nlNni7CRcxN+7CrD8OvGgh0lk6MYzjESKG6IHEC2qxYp
0IzbvYL3SwWfial+Rw25p+Tz9kBVvm6JSnwDzvthP8/CriHrcPQ1SJa8jzja/lLM
Rh9Lnq7bKJby+Yj9cG62atEfsbLXIeHIbndMxaAJLNyeWMJhhPc4EKqKB/UoRZ6V
LTmITj4izwD7IEcBPOUZ2xfz84AjA13a12laxkjGJdW9ICMxrvYq45M+QkGxDeqZ
KpQv1uQalCH/WeXNW+dAIytMKs7/fWyaqd/SMn/3yUxkVyid2U1HL2CTFj3imNH3
cCHrgq6zNhqL+rmMZq2OrzVNNpuh1biljz57gtdPmc2AxEfdB5X98v+0ygZ1Ec/E
laOeHdetqPPj4Jv/xa0888pjok88FDnjTX1uCi1atMHtEZhdbwTqYVzG3vN98r38
6QHEiqP820q2pwbPSbn980xgpnYeRqMg2QFW5zh1XO9bK+D9eG3e60vVfEjDD+A0
mNhIuKInxvhNSDcNMSnv9FbREh45QTSOastIQ4hZB79YUbTIqygILM5x93OcMoHs
Tj3+RiXN8TxESwKNJErdaMyzb6QByjH0gZFvoeKAKp2cyB45gzf0imPP3HUJ6wU1
jC1jU7CWRNEP4CU70C/HYPAPTLjzt6B0tYv+eJMi6nHHaGgn3qdJz5OKDKDxdzDR
+h5PP0X5xYSmx6HIX8cDIvvuk7UNc1YF3QHzJyV7xOb8rMhcJ8Hb1Z+rTWv0+PHs
/Y446cm4kGzkyW91+6C+Cpx7x21+lJHyZ6BK8bPFwbvUle1b551j32pDPSsSJO4+
VMkDeuzShwfQDZvy+DqZ8pcrQfcOse8bVKIxkitMkqYM4G5aF7QKDUZy45nhP7XZ
zPwKaCYxmAz4edLg7FokwQQJYHSbsJdw62HnNt2E9VUSfiHaxY45EkzaxW+1BY3W
gdsksO/Q1vYP/uwpdefbAVbCYNf12iFfGP7rCZSadWYCT5Yl9uhXCnBYtlryBULE
hwARZA1H/wh/0H3NyNobz9oTTFavNVrgMWf+1LCWVU7bP+fEvdqA5JWBv69gnPSO
2qdx3UnBX2peDTWJZ2UQFEELQEud6S883dUN3nB/MCQdiFbITyeqqZ8FCZY+HR7c
QTIVFJPBx3qtB7ULpy4Iy3t6bT0YYONpznro7MoCMYN6VCZTSK+D7fmVBk8H/NEu
yko4q3BZzYFQ+rQ5B4T3+rKn5ekbGVoAP1aGfePLcek+ZPJFJFwg3FkQanUKNzPv
1DxZTL1NO6eMo3E6eeauS9akxy93IHBI2hAdZxXUuIX1I5RbkN8DoC4U9fV/Pr+p
7wp/+UAFGLfe1H9+z6Nq4u82r1n3lNFj64QZu9/1wny1XS1/u9ecQXNytVVg0ald
ayWCGUDZ1IZBsa59hRQG99SIiICw/teh/Lx2txdT8S4dzTQWqPhz2Se7uUT1I+1w
3rXYRWF3zG+V9of/Jdg88biMT6Tfooli51BrJ5faxVjAsTz531uMpwgh/mlONgbd
8zYqcjwSVZkCEUKemr696axAO1ruBMSalLfRiObiucShHOde3SGPaIAH3mT3QmiP
s7biq6BU/AeWCNexclMFGCyiptkYT1+SgGvT8I1ZDmgPCGVlxzU9y4GZCHy4bttL
82JjTEvxLGbj6GYPtWlSEHMBb9qe5hW7NyAZ+jA9pWBC62fUqltDCOi4yHv4R+Qd
gzVjMlIPOGdeZXsGJXT8eYkmNLME+ZxRtG8ifKnJBh60PiZW+7GdAa9GsjRGhwnB
9fHamBW0RV9DlQ0x/fSZORCvZxxF/S9LZTqaAgBn2n/WRMt1jSkT/+9kZ8YF5uJB
NiAv32VENuz9Ax+zeyEOGPHU7zb56KvJ/yZNHkqj7ZP19MrKibgQRm66dln1NeIC
CBAQLt67RQ64eWHZ08U3+A26aa+6P4Rew5FFQfiqwogkfGEyz8Jz3lw7aR9dRDg/
/2ez0yXesFoBBf9wY17/Gatsxjhf/dA3lW+/EhmngwdEORTJyD0WggFl1Lb9z9VM
B3zaZGenD9V0514EFTI71OkkcWEHEaIClEfX3nMlzjzNYfKNNKjNMOE8qJvWblXc
InpudNK8+e7srUtiwCsm8J3HGDBl/5KNyIWNcvaS1Q0mA2vWZn4me8qKyj2uZJwn
di/J7uemllsjSPPc9ss5gBJvlfumhKrnYsTdIS+dVtx9/aWWRT0TgS0ykSukr51R
Y97zgwkS/W/KKkfNaZxGcuntdLgoObgrYNBUtgyghYiXL1dAVo0v1uGkHSXDV5Nz
L5WipeR7fpneG65FkQOjJeoAuEuZEGhCDo9Bmh7mg2zB9OsdGRe1+Mm4CxNHT4xG
T0XZF7ChcRx9yCUJaKrPIbQT2PwMbwqaRMzsPBvOf9eTqsuqrM9Nn6r+5OOIpEQs
BmtLoGwsitWSKnWIGlfuIxD7hHA8CkjYAwTG9Zada49x0mbdWmBGM6H8HcYReTMG
tdsDMPxV175SqbuSo9G0AQz+uv1cKEj0keYqY8Y/oihNMe5ASE3ric1XCJpolON9
E34BXsx0O1jARBbF9BV23wDFT3vHyrUa/BMENLNSSCNOYFr/myERL5dzf1lfXJJl
2D7Rmjqn73hg/rm0HxUCQD6a2M/8Ono6yAg+pg6PD5P5zC+oxfoD0NuJd+GLDHcU
I1JFZgXkQg/Rv5RKqwuVdLKuMCgowiuForIc3St66lg64q0kzoheZbRYoKDTcgHQ
OGqJcEYUz3spzJzdwFAQB0lTbGWAS0PfNvIpRuOD7fk2bb+dRK5iL5kw9zeQWEMV
P8eh0odFbRhKwFPQF5GJQDcfqtR2jpSOU4fiaXeivWSsiX0mIkr3a5/vSUhRi1OZ
JH2qORmRij5lMMljXQZ/9p4UTE3k/5NR4Misp82w0MOzH9A36fx0E05HRZzGUmMS
y/mKKcbeQ5y7rhtnO4XXi2siskBs+5AV4YYlhzZ6E9zMw8XerEmTV8/+sOauBdli
9wg/jlH7YmKi0ZnGdfnAbJLsbGF9qxXYyi8bW+39r/H0p7Op4l6eoNldCYv0jO6H
XlB89MXx//ftXbsQ0HZugVcfPe3clM7ZbWf1mcIgOK/+rJ2mSgcO79M9ajEP2M8Q
mZKEoUYOJT7bA21ofZz3YHKj5l4DbqyUFc1R6rxK5IdbqfIJAKvGg6Up1IKXT2uq
vqWibZd7nMYtvr/rBZqy2DA+T/RESN/a1Fcvz8HP3W1kq7ssxLuQ8Ezt2S1zXR9Z
XgdX0/r+vjuCy88HzYn7CZaSQLz6XamR+V1wW+NJbnbzAwA5QpL9xKxk5koztPkZ
96q4jR9NtLqedYDE7YF8tv6RizeEUdALYEKifLPmeQR85cszC6YVbu7JduXHXTgn
oeCJ+NpwUf7zMph0cS8brPnuPSG8isK+9NeBgg0NgmRGgE+2qjxgqtWU4y2vDwob
P5rtL3aMUgSO/A78R4pbvGgKCHXzLR+mU4H3+XwdqEOXkqKmdLrPA2vAHSvICIG/
+KKqHtFHIajBXpsFZmQ3SLpLxAadx/TZ2AlF5vPDAtBW9GvEsHzFo4s0a5oo5o/t
hVQhwSDgRr5+vDwL1fwhjHOHtOL/v7kTr84g2w/KJg6gI9HbA31e3IbZdNhAolxl
MGmJHkGqcu7xITAPQ+Z4a/GbF5btA0FDZVaneYa8n9gxhDvSAsmlrbH3ZQmxAnpI
sOWDXtbdFg6ndNIsvz7reCUK+/K9+6p8RqVLJX2SAPkATbRI+NfVro8oGJHjcveV
aiaurKzz1+az2/JSSHWTOSgJGXsY27Qob9V/XKWw/5rLY3dGTxqlx6dRabBgqCjF
o/7OMl1uZPKr1gV5FuAXTShT/dmoktnogNUw/RqisxdephIJQL2na+zOUm1qC+Ty
atl5wZWaUpuaPEGMdocj12ieL2LKoy3IRafGHDOqolLtd0Brp7Slm4lVqOb3mcvf
zAilqlfiCErw3Au8t4djV5aDN2ZY0lIsIOBDpGjUTmRq0lAfcrNYQHpjBXubjdbh
yQBeptJX3iY50XcyNR0lAeOYpp2k5g3HmQCisnplDuW5PuX11LdBY4lGAzdHO0B1
89hzTYQEV/SCRvpdsFz2Ex80UQe4rlHDRmohxn2ObQHQOb1nsCtGXIDeUO3scnVM
`pragma protect end_protected
