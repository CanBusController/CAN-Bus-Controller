// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
AH40OkFJrO7Q0hpIABVpPcRaERilsFd5T2KPs0XvS8NITmRazlTFgMDDNKHOkZHqNDW7XU20YhpR
ids1NUe9HcMmT/8MpTVxULyFu6UTFzSnH+G0VEf3UNPpwdAJHH4xZ37SXNJGmiTm1ImWQiXc0/A4
kcfJWFrKnNA1FTfRzP7/TwA0veNOk0+6qW8WpbPIqF/z1gqy0lTY776BYx8xKwL7hfJ5k8UL0AGO
wxQXAQI68yLn3j/ccEnxYV4524PzQv5sgPexi7H9Z1It/1woJ1mf7YuKFwkRGq6W4ZRxMk48pZvY
T3/FO9WzWJSbZpXdW+EBifY1EDOmwCRwgJbHiw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
5fIgH3X5LrrH580PgmbXopAfhzOW+Ios/YsI6NuDTQxcjBjx6BpQOGCRo4cNap8zqcdpAyiwgOsM
mDhls1HWeM3S+LI1gQBQe6f5kGBDkqLn5Z7gPBXHYfhvjrqczjA3hFdahN5viW9ct9vv1Mny1Tkr
HBwhwAkhxy5Du6WHfPywn8anygwEHDfX6noSdVYlrXC7W0HRprlnAShJbtyF84w+IcTdOtfUxwyr
W04Pl8iYEDJv2SyOCBciFrKAqX5dYqdMh3Z/AKT+93eYUTahdbL43fXTEjSkMrU36vcMprSy36uL
dYejlGGjVa8Z8oqSB9WYvBROJV2sAH7Oebg3FdLeBH/EdRuO9NZZjWIvZ0a88meAgUjGNaM4RxPH
SI5/+Y1txrbV6fEtDLwv4U+woQnUM55pNtLvTVWpzyaJBbpXczqepcNnUKCadJaZuqhLgm4xORZe
wRGLiNxa7p4MjNDCVmPPirdH0Ru8uEEwFozvO8p1qnXL48w4Iw4RGzhqYJYp7K14rXYHMhdLGbEb
ID6Z4JTE6GFNvW7Rrv+vRFgCe+wtOVF2Vp35oJaQBc9YtD2stWJK9AHrj/77aqr8jpbZ2cx+B61N
aksSiOxPKEQDm7glocCepdY+9cQUP+9GHzpIP0+aZ+Uj546eLiav0uKIKq0UBIfNWlMgKVtUpTLO
+Z+EOHz6mxnmSu+RuOkFU2pMCp3jX0F/KwemtciZuSRrVEIff8bfG4LObkizOCU7BV3kgg4lBzr4
QjOanBB8lkMK0cXq1rKHJB+knp2THVvQzs9LcBdoT3cVh0P+t4D+yEsLjhum8pRn/pQQNEnkwCPQ
7vH/AkFiS20ht8MDomDcnunQB2+RTVsXQKwU1AVjDWXjazMjLz9ARs7MhRnifq/hUpNUTUiLwg8J
sD3cuBD+ouueIYBv93XqcIs7yz8Cp8LXGRDlW2Z8oSX7jOPVCmOcggbm/3tGPI1V4LOgTKjFwQIu
rHCajD8RNDnXEZMwrFL6I+gr/+ynYp8WiZXPGTyQqt+1muFCBlLgggOiBtR3ZXAchMA9qkj7Q0FX
2BSJMFS3mU6OQNrmWg5yPLcfqMV32VchyX6AoZ3gAZLftYUGuUiNAk34/AOaxbh0L0baZefRb+ga
ZV0YJsOFDqOt7DxGmgxadv35jYqOqHXm9kO609SrGSEnMDWRIHpyZKIhMyC1+S1SL72BMaJ7Kw1v
t79MHFpoR4D01Gjwq7MqDEBcAb2ioR0rMI/30lM66gy+x8IZ1hHlSlFVDcnhg0UtzJ8qPNIf1jWY
+T7ytQcC5XZIFWI8qN5QT58PenM1ZVuPB0+MuBiymFqPAG+HMlpM72Iw7KopPp0kJs8Gzsna+IB+
di6P/QpyGg/8nwkrN9bQldVq4mCw2vJW6vj94hSvv4AUSdftp3mi4RGtDDAWBKGbjnt0U5h6jNFr
jwL6tModwII9eoXgQfklGVT3p5n6lPHNLkEDu732fLxHC6mSZ4tIN7CWBFlTWfjcD1v+52q6gyoA
jIrsBJ37BGHvXkTC/We+OE1JDjMUPJzMsoWpGvD5tAzmaFdsIUiOntktHcZGHdgQBLWbQsUu2+zO
oS0S+AKsx4b8QynX4NeWaVZRy/UiBK0WSbPBQoOL0tsgdu/XBm5wfRiibo5TiMLwzhdF/dAsVpO/
EcNNrIfBemsogdlrXhmMkcW0W1Qvw+eDyoPUPPPuZVClDrRx4gLvWQF+eje1/oe/7OsbOFD/CIk4
BpyG7WaSNBazBtI7csZtDwRjRTJ2StYBB+5+ulbzQSivOf5Tqpiev04DKNYPuU4ors+HDYuum8o/
aMCn9g7qcl2H3wxbNly4O24gA7/MVz9Fj6wI/DymB6V5s6Qitoa9SJsI1vETjsOvlXs8aAa1sIrj
DpiCN7YMF9HPsd6R3RrBKROW+kxuT+ae7n0oIKWrHtaJ0oGc64GGiX52lMK/nHmpVZ7bQfK2XSkO
FOFm2ZoqSXvIg4M8HLj8t1cVaayrN4NbGq3TM2wFrWaphHSJva9f6uqsLF0Zq/hlyuNrAHMiXWkW
3r1JOqPR1nh7SKPVxgT2pPQYZqN6gwdoKci0v9qNZPCTqz48CpLrTaGdGL5Kl0sQGHUydcPFLOm2
NMhM5KEZfZl7pNahgUhpxjZUH1HhjFAJdFLMnU2+Ouu9U/7JegX0G+tZ3jRovqrLEOC+z0J+0uDs
U5SRkzlQ14xr61nodojw6zXbz6SK9M721uK1Jwv9s0z/M1fOb2SlhXTo80wjEhm9wOdPan79FUJj
gBuoqC23stQ9zrhkaF0Qw2DrUYBfgOMbj//CdiVCs31WIgMCBVX83vun8JkXfXOa/8RdMrxLE6ar
+PlfBDMHJ4ZoX9Kxcuk1hu6lnwMl5S3BS8CG3VJ5MGkpdZcoPmkSNVpYUJlQmwweX0tefXl7Is0C
aEF7NeVHRSsnpbb75/jQ+N0fW03rlKE32MvkFj0+qhDOgxCJi2PDFNA0BiomUTyHEMjfazaC6tzO
/0RiWKpcNDGe8oGNFe5u6/RbiLaNKUv2Rh6KRLBrRDTwOoqn5ehVTHAY5TvTnglVJETQzrkN3+b9
Arm8O7CovPCdSpb8F6NORS4BnJX1x1gGbRtxduaVt69Ve/s/gXcoxfbmmY9APmCXa9eh2xGQXOGJ
w4/VnqF+KD1jymsj+zEm3jwLQr+aQrr2Tzg//yRRbWggbjc9pHvjxSLI4tbpNtRzAFeANzgS/GYA
vu2gRpdL+uanARF2x86GSBzBvPqIQ8c3ZX9i24rasD8I1MqdVa7zG/94PP3ePPnEmTODC2G/U/tc
KezPp52oRLwBrHMCiF1dS8GZW61V0oMfayaGeB2VTtI4Wh9htxfd4dAxp5DsrolXMJGnqHY1rzZG
YPZvpmLT+Vm4Ts08UGB4YUP2OlAykhSM7dd4BWwpTpn5LCMEyVSM8BpcJ77I/tXBlHK3Ax/wFI/L
N4VeEiZGkjV9qAZhgXqYEtGgM+M6tEYn2x5JJxTkN3R5VTn2FyzbOWAPBc9mSMPyn9YNOBoXyrJJ
nd4J49QtSfXdrW3MkLGU5A1ornpLYA0/y0BFceem3KpAN29mZpTXD5cpl+bOQAI43Yy7MQjERxIw
ekOakWwZ7yYdnar+B3CkOZUIe/xJQ4g6s9bBNTVKnu92VWePwfw3ZsbY3qrNuw1jFeP4UVHzvtJK
nclQZcK3njKSti9rXCPJgKRHYOxin+UWHqaaUx4PP8W89rk/uJtlCUUnjmVgnyHCPKNfp9w6/pJT
ZGMukKhbCJboWEyX+cljYeU7u7XLMXMS3n4oDwl+9HSQHlufAdjX1APH9kIUHia49/dGEbpi/2X9
kfxCE4wZ2pHBQmmJ5pJxBsIlit2kH0TDhA5dy0toml8g/wP4doWnfWzaXwsLkChX25LWbSGv+FCB
QVSXYAMnAjrXMprZGqvItlozEofmH/8ZDnoDE11JV4LN6TsFtNe9TUZQWDTKY55MuIRuRrlIBczp
k+XNNPOivdIBt0F4uRdW74Y9mlJdlgqptiR56K14UcofitN8tQr6GAz1P/gmiOOu9nJn1X9WpzTG
VGtJTGaj86yVM5kEz3UQDRom/2sNU/dn4/gzWVOtcIGuyqva28xPt9QoqbPWXgiObUuQEP0G77BH
cdM2owufyIJjI22hN16FSe27boWIcad8vf4mCO6SMu3BfsnMzb/EhuVnqhBByJOVQiV268n6blt2
MwNpNxcoZMBJ+Ur1O8IawHuieFj6uWlw6Da+s+oU5RDg6+/S2UB3zmibqViXmC5zn386Vp7xGQtp
4QHU8F33dkA39wciRM4KF9ZHEQOWB3qXAmz3lztDgOdH4m0n7pPEP5ZUZHcT/Qh/9cxiezVt3ZLP
wLjz87eq5/QvxpIzAGdrnLuGeMV85t8wOvrJrB1v7x8zGm7n29HlLoLIX0AsdTYMVRg7uIs1JBCq
EuKCayzUdOMft4Xd6i0+Fodl7rUSMoN2t9pafqcyd/OkMDdU7FvrRF+vkD375F1IwUdgjv9G2kP+
iWq+LTgW6stxuwK2MhHiVhW/DFLbrNI+z0NUViDrwNLDiryziCoPXto2+oVxApFxWqC/I9EVvkqR
gNs0icZCR0fDvoMrJcm2g5XbeFUhOA73q3aZsAa5ktfK/WUgpm35wQIa1zqYqXw9kr1OjLsiqXLr
87ss8oK1djHhuETRx2ZBSo6gj2nuItffJbKD38htRIlB96MIalqN+H0i4+trPb6lI2PFCivuUqxS
vS1/OQUnemgrlXmD67sc2ZxVtQ/fk4FvZcjov8E5kF9gklPH7Ad7tb6lbIgsI77orcuV/2WN7ytG
VJPfMnOCoPwZefci4l62k32aklkcxVLGLjE/Tv4TSPm0HAmBycKnKDzgrs9axeE0d/22AAwLi3Me
umOxpjwkzl/+hz1LcW++MhSWjtwZ8meGugzJEO6aPDTzsbfeOPyYPsKBq2cIVbFatG+2er3o1fbZ
kreWzB331cR/j3OO6d6fWoqMCqRbC8/x0wavF2ERo4GuGdAQBxeQELQgO77abm5H9e1rLRNMGQ6Y
v0jGTl4p+w1TIomEOzIx8cbFMxPsjldAKimnkmEbuxOpC6201GaXdsfxZDsFBOjL0GGqpDdqijso
doQtv2+ug1BkaOUXhjjPS/jWoCIUq4bVZ+NfAscbdKCDUpgbGjgdCUKfaJo4MntPDzG+zZExV4pF
h2yvhKhRzNGQ30NXgWcuqpVhnuyR1L7UyeH7NYe+a5qrCzfpB1K6t3jGXYmRrLBL1xfX6TcoKBPl
WyB2gGJbPrxoZ3u3BabyO6qeVbhC3/ZielqVwKnn+YWmgxqK6yVXTY5tVX3ejoNdAHznvs75IrxU
me9WHQUYjYuzxCTE9wrgKvNugGSB9mFm+HLyaqhErV3xaDe6FxQB4c0BxNfV6q40SvWIA8WAr9+C
dToaw3Woq0yHNrb9dasTmD5Uq9nnJMh8uX49ZKWWbXp0PqU8QaeuISHVP7D3TsZ0f4nLO6Ry0IPn
B7wpN7LaF9+1YC4/0Wv4H+xKhN3xn1qTuCrQZHgjeW2yebTfpPFU+tIxbkAfkufNvHdvuzXkxXqh
D/64f5CU2fIoyix4ouG3oRtM0/m5PL25Wh8nzOvxISjRRpfJW8TygK+BvRfJ2mQlgcgc8qy47TkT
ja9640JQOHrxI7/eG5GvSvBmURBnorg0v/TfWVeVpcN0I5S5pqEnNhhR5C1rlNjvv8xHJIXfr5y1
9zOJ7iknnTL0ZfAGmwIPzACsODVuLVfOuYRAK5Sko9L61mPdW0S7g4VWXTyD6/pqkRqVgRbgz9Xa
srDPwjphc8O7FW4F+nAwZGTRVZGYN4aykasQR9HnN8V/aDkI9XfKx6FMV7YQrwtKtqCTa8IttbsP
xQM7RLPuXk/qXZRlgprWTJ9wXRw8VbiWIu8jLv5QrnNixE+JIl9/eNq3SlEq00jdU07audB+DtCf
sh73Jwln0w3xW0WlbiuFr0oRHBkKBSrGDpjs5NS5D3WMRlR4fYpbu7tOBR51nnYTiHYF7a/ntLVt
Wwn4YN44ao9+V9cqkFCKz12kWy6WXxXmzGtTvoJ7ez2CohDyw1DyB7jTnoJ/Q0qcGrEMMCBQapEz
kJFBX7/SE0SAP1mmVGaVdF8pH5Av6gSQzEllVifS9QikMBy1ll+v6WSnXGo0UDhOfX71Veolloq1
dCgSfPk8WX8F4P+vggUeE8xKnJCb4XejGqd8Fy3sztM0+mhnH2skZMgwLilYIcmrhHNoPc47o50p
Qu34vWe/UGj7BvULHXBu9NUjk4ePkSJJNoa3ZFKuoZloIFN300B2k/FYDzVwyqwGuemqLolSV4M4
QgYpn3y3hru3+yPAGcztaOYBGoBAKX/BEIikhW0zzLZ0nYUhBRIBLVzY2FMaTlpkVerO23INm5ni
EZU2onVmpyvCsWTbNSO+CvmH3QxWO2PofPqKPSoHKSoYSs7PgSR/XRUTNmHvNWmZXc5xH+vbVguV
nHH2d7oa6qM43uTspgLjcwFJgfqba0naiOejQSMOJcHj/4zc5aNVFsL9Ql20nHVrZRo++M5RDoXz
AXt5icjsi4F17aHkWg5BaEMucZR1Fk+03UdQ4KFPtM+iS2AB2FWo/WbzJVc8ChbKnx9ZNASKTPU+
X2l/LzwLqWaL4DptGSAPKXz3rE5oPNwfguF/+jvA0zxz66TJDjXd0DYfWgvHHCOmwT5HCLapYGy0
7dd4mTelIxUpdpx+4+PFgYzG6egUIQkg/TiB/1PPN0yW/Rzu18UR886CWzGZpaEnw3aJsJ+YBxNZ
dt+QbBsJIy9TYlq/MMTlHJzC76OqIW1E+qpdgtQm5OBgotD5l1n35z/ULoF6xC2HiOqti1EhfI78
9FCRFD63sRppCDE2H3LWrPYcRPB6eLuWdTQcUCB8iVf+NNxaH57xcvJ3Y5LfIqbW3WsWd+8Uxqs4
7bZKT1L2VWWJO49oo5i4l5xx2tHEaOLNSiRpwa/pGhm5/a2XFuBvI84+uRx4cIZMZw/LWq2d3qn2
SJSzaH0sQxnOFkuBPPGQjGgCnB9Wnr6ADnUgDcPuzy9BAljD0ROxzXWZjSYhf6R73gVy6eXJKMeo
fG1e5PVvpYLBXUXbesmg9jQPyWA3uikqkhr5VWtJ6TDuPk8sFNE5rMp1C+olTF2gbhcx0gfLyue7
MIujttyXdGe9rWb9NPAbmjEkD2uySe4IpomKsjEshhFRdswVrcOCzYDXBoE0RFM69h/fT5ddPbXv
LpzRGePR5yvt1ctV4ED/o+7l7eTambSexyMIihER4VLBqFhG4iSKv/mHheHN40lV1m5VfJbBZBpV
0OVPwqVYySSfYGR1csqsMZ0q2/jGawl/CyzWF1fKEh3XafVAAXXs2Dxh/mSFtQZAWlG5JjNaQaR9
dMrhVqMb+wJr3KAomn4w4YkSla0XyD4u2YWAh82oHKF1jzFSDXJAK/EgC+4YBP/N5wDhWHWE0aTm
dDnUQvHfb9Z0YMyKCKf+W05+JdMw+a1QpV6kCDssdrhRatTsxzNiiIEMfv3zf5E6P79OOEALLjRD
XaTFseWbRRo2i0SdwdIo+RDCoxcAaNawCNgXR263nzqxNg+RxZU67PxuUWph0pSoDFQ/plHXptOx
h0CPv5v5I3R5PMl9g0+xfKjS/VRJIWA9cbSOpe0QwKRCstv3ev2QhIxA4Dm9NHgSxMS8BszLgg1F
UVX3xzCQstyLOCEmdi8MWwzJIuqj6RYr2WoBzIcYKhhfdWssS4v94NJzJiTSLKWh5awFVfd8ZMTG
EbF7MeGCBvLmxomT5KlMYw2N2icmWfzYrGfrnZuhQIBzsSKfvKtjSbSg+XO282P0o1XXYD3uJMiw
6xpIEOz+C6JwAVxeNdqVCT0CDJkaaNtVp/gNtxHlAdTcLvxtoQqmRi1J/nhM8OZXKGJVZ96tOHss
/DWbLwFfV/m+3EgHZ9UtfxWn7ceHVYziJWIRHUYmHOWStiAuEeQ941Z7tJYs6cXftIqUTdr6vydQ
Y9oY5O3JKlq3pFJn/z/8+6Ywv6G1aTpBuVcZq4NANwk5oHFVQd4xo2aKh4zCKZVmQmJy32E53kob
r+tkVlezrEokeYaS9E+VU4D2bcIWl8HvkNxktcn+KhFEsSLPG05abLUgkyTb4SbmfmvBu6md+ObB
CapKFoQYlh4Yq/wSJ/G9o7h1xhcC8wqnWd5HpBOmXB06qbBeEEOJaN0HT/7QoEzYWBkTctqeeeN5
JYNx2aGjaSSS/tNs9K/vCL95koIOd3A+KrzH8BlyxJwgNTVLpaw5YhZBs4QP1Tz5esRDIUQRs2Ws
W78RTQ+mSZxdSWRnxkdYPlXHB6aoSAkAUnAiosG6IEeCXFpH80UVQ2ZMVPwIUn0TosOme8jRmwmA
v+aW/nhZc/mwVKuM6Zu4U3MKsCjKCHk10j0pIiuOJ8wHAfjIFdkEVBd2yR1dSIjC/mL1sfCYcIO8
kdMrj2YACTu9Hp1FzbfMY7kwSFfntlx1ZAtTfYtkUVvE/Wkv5BCPT9XXHJvbR/M9RmvJFSgIsuLB
vv7UexvbMSMn03vNkrKtyEXoaD9pMhiok5K7rc7eNg2fFN4lw6Ug07K1zklMulMx9XUDxcX7c/VS
3l0xIVqd779ZbknlqrZ0XYVkQIvaKjYAM4fQSE0E5yMUFua3ABXPCTAEeAGirARmopoQ6dglU5vJ
vLN3knM17SvYDe0sOAgNs69ABwtCaVHLRmRVboFdDE0jzQnGJqE8CG9U/rflIsMjhJdJEpWduY8i
Wrr7zjFqyfozcVkJRserbKm1Z2jQ/weRBlfZ3abUzGmVorysULfELjVLJoHsCdVZKJq28zSkCjRw
9Zbsg4Cg1o3Yj9b584QJ4ym5CU5ngo6TsLeQlzJR03JEGeqc+Kvy5V45eF66WNt7mCvRF35yqtgo
WX3MauumaUQz+DdYLbvUajJJRv3BO2tBhI33dsI52CGllrQ8BaqZDqAdpJxxquin5eTbH7gFD4d6
Zfxjj93Q0WzlE5GsOAlLOhPYZvvQeC3MLz4dPFOy/Ws4x4eoTS6YmdaZJJgLOF2KeuUHfEHNjFxK
1AtrpYATqbqsR6MCiFnefY20ZIUKEBygzP6hG6V76hBl/XT8Ccj7cz/YCOrHOpyXq0Dev3c4aweM
poCnb/dbb7XGIIvbdqWPx8N30yjZgRVURVRVI1sqi89mOvFD+eDu/8KCdcPnPgEgxZ7+ADfoy5Co
ihkET+9GnyQrnvevXVtoHcSYG2qDjtEKO3uSBtBlphVWa2Au6/QDN25p4k3RyFJXsS55bpcgSuVb
N9Y8cwncFzREsz6ub/Q420SzO1Yia7kQmWMu54aJ0YPibONq8spprhZ9SYYMIaccSB17Ffga2ciy
QmyBq7H0vVzAAgH3Cq91CKGQhpyEsrk3YUa4xDLX5z74/Omvb29MDT/uIK+E5QfwGfL5rIyR/kM0
cilXEaZcvLKlBAvJN/TSgacuWqBTfc3AoXVUUI7VCkm6DR2ZuEh84QRcFPXNK0UJB48mNsT3mHdL
+LmCYacArCHtOeGXgjRBNtTtwfZhc3uXkZYXWe/fRYY9wl0tfsni6VDTYnkskUcPvllHSLQ8uMKo
pXlYQtjVK2AzO3+3ikSJQRCe7S595WYOOPOXsy2qy4/z8iDoW6Dp9/Rye0qQ3nnsYv6fNfqZYmAK
1EXYxxYwKqnHRl6NntMl9r1YwWyG9KI7G6v8r6AtdSdKzYO2AdbGXS+LqtAO0f4gGo2XEr37oXMn
cPacWi1JXPqtPBc78kkcL/vbYjVN6WiMtmizn+UWmNz6YmpOWBOSHn/cnu4+PR7G8GqFgf/ZbO4S
hep6dr9b/lHJs26z5jESB3BG5ZTERvgMXlpNGEwz+gl8ovzqJ1/87PE3SVetqIBV60XKSFhbTYS2
4zaO8MwgzDJlg+NO4VLWQvh2wqm75yucl6fHaemnjvWV+INCSw4ubuGhcLAFF1I3eeVl0IQToYOV
BrjkfNIImJorqjYhlqjdSg5+Q+1HMRvBTl3onwd7sZzwzkDPrb5RSYScsPfdFZ1QbcPe0gk3sb52
PfWaIOg4wcU6GAE/qyhgfZ0Njh0OCbrUSuY8QfvSOEIsrt+ehPoH03FhxVRXHHnOPmxtmYTQ7wzQ
aj9SLnXImKg2Q6Bf9xNPtFchbP/PAG+oAHIy15/KUQLFuX0Yq2W0Y7Df4ao/a9ItT10DdFSuYvOa
Fri1DLpVnrwNYMHPQX8ZfY8RwUiGlsRloNgqf6KWI7V5y5gWFmN0Qz61cB04Ij7dhr3//6yVAOKG
wU84MHjPsn4eTYiYUARt6d7+k7wONALRuSaj2/3Z7K5xaqujWYqQ75dji92YBYqxevd5FkHB9BEs
rIJLLbn3OGs94U0oX3hB8R81xI9dM0AkRoxxjAgCEHZY3wdFi4leLnZeTMdNIq4124P+kxSd3wmD
Op0DQhmWL+ROpnoTIkIFIOlOoa7MNLwfeRs6+XP/OIMBw5LB3MfXpaICmEDo1NXgQz19/YAHWMIc
J9fSqDmztwfSqiOf5hEPl3pT9Lf3ZFwl8SpOkQsZY+apSBlZpeqyV+n1qtUA6MoumyabtBIFx2xp
3xIrwzMMnQN/uCkMsL9SmSNUw/TwBLgWH5y60tqI1EyoyMtfMkpaaGmdUsBXMJ7AvIYy/Pkv4zVp
smvHbF/VwPKlzHqzq/BcEFOZGOhjjFnNWZsy+EU6mG4lbelC48W5hpDiAr12cs3Epso3bJIf3He5
l7sLOQj5wWDIxGLe5i7H8er6IU1HPKHYTVAygnXZ8a738FZ6gk0xLrqdFnyW//FbwK0GI4tNJ7uj
ggLCqHaK5YtPw/txAX1gdlRUvMQs+NVAt8G+EAD+0kBUNJO1vSheGUvJH07m6mFbb7isrkBSBl+N
5PLy4UGxBWEqnJANE3hO3iZuSaSLbO41zh+Q0BIUCVbN0xibEGdsCnT8PXvirOjZttoX0pCdFPA7
Zc3vU22K6S/meva0B9f3/lSMMBOkQKGJ4aVsOE1WuNUkXBmHqAnnceQCYShy6iAqpoodPOOugGpc
XWWw4duuH1Mfzmeoks2GCMj6UsUt7oA5rvOxWo4ht2g2OHg9d+ZuFKk36QuVP9ibzPIqpECrPorx
GXTaQK7pP1v+D1iIZR1ZqB8r8bwaNqR3ri7e6bPcapukkJJ2yy2bXPUZLSalZfT4lszubYn2uVAA
2LzWVg7HMA8R1AzDlPOwB1R/QkVEWGbfo1FqACHiXb17QAGEHseMlq+WTouX+whfyACPwqTd0f/7
tsUxcgtEvOsIDENXVn4JYSft+HlUN71Dl9H7GxEDQEf+ii3PGv2+56RKUsnvgzjZ8aRSe0FY7v7A
85S9aQrdva6Pjxa4kNfhTDHz6/8LCWgKUY8k9L3AWBQNv1J2LEALfkrWSrhb4p6X2jVCqxYwPddU
tikXntYSnVr56+sXYUAgctVIYJ2/qYtwwQWx4xd21BbbXs3mZSN/ZkBuc5y51L70ZpYqdbd7EOaR
pPOzpunIfA33bFip9eD1W/IGJuHKME3SvN8is38nYq+bK/W1a+JR0LixIn/A/oOXYfblYgKXspkX
RGjLv4wsQKia3LEl011Fj7b626sGL8eOJQyavw5T0UIG3BVi86Ke3/MWC1c87lDcask0N/AIxKMe
/RgpUItWrzU/szESy28tleb+xt3Ju3ZodzibHpF/SnxX7kxQt4KrVzMyX2n9MoTtPNcZaMJ69oOU
oQYEzMMX7cgNUN6ZPvTqZbFAZ+PG7JYgKqDofRG+VrIqcfHYX10SUdspUGfbKmah9xT9mRChPcc5
mArJyb+XUZ87l7UXgDJDLMQ4JKACghijeFfntfUkGEu8rpPfw52xoJd9C7pgLgQ6cF3PJkdyAD7+
o8TvCNR4oD7grGsVTo67wwAHJ0ze3zncRY4Di4gd8WaVmg1fOe6o31UpCG451GgAcNfAbZiiSMTc
QzbJtDywyWTfKp7D94FcDwNtT0WdEhzRtlZOP6RPX1nKpvjPvy499owntBoNGb7sQnXH0owvAQ+g
qcRNs9nazolo/EjuCl95+9YTRFr6h9e/yDtvvAT0G9BXoHCMqZ2+vYyQFnxHty4GWQnnn4s4Cgy7
uz+0mq7y+uEXTdrew3ewAfEYCV5/Xebi6jtf9iKj5TA0fSt0+M/2Pj4kUVQrHrt3BXxAKN/oY3Wp
AalKTsI3lcaU/uTekm9S2nptcNKtFiCwEDi7E86/UKG7b3FYAFWvDZoO24I3BhKszTCmLomiblDc
5rthxEwvjXSPBjKhXAkbr4xiPBMglQfO02LEgVrgawVdpQGXSuQ6yzMyEX5tdlgJpgUAGW7h9qsD
h90P0dG7CrpkySaZ/Opvb2vh1OHmsUdTVO5dsZ+t1Qd925dQlGJnsXYYvT7eV84stvpNzktEwYr2
xRYa9pXy47ZUuX+Jeb47MpMsiEXGOZLl5DIQKm60auq5L6I44S+rIQawEx3XJrvKTUuHgW4p+Phn
/PPZfWr/+fJxACAhwi0ybEY88dhgyWHM87l6s0Aki19uiYxUfHzYPk+yktAnSN/6+Fc6YWtgKlok
ISRmh5xJROHT+XfVg05KWoNaPhAXHBNR+2MhaE//eBl6VtQAs+752TLj56KMOxhi81GszEz/eL+T
AxEXb5aD7S7lQfvfQTOgw/TOWMhCVbqB66gvqZl5uDmcH9Gy/D2TRXMw3uy6O8Zhnu2CA10bkYrU
ihsDhh9RQMlqoogLnPbj6erzuSuKjKDmd23oSwKQwWygLGqOf2OZsCXITLcn6q3EZ7L8XEw7VW6k
tvyv9Mr6BLrO4poqrfUfK7zAehB5GeUhfzXWSALfKskz32kqqa4yXBrV38Atd4f7Z31Bq8rux1fh
3ytEy0WS3dPfpse3JpaE81hzOILILyeziPEm5lXvrIwgevyWYrBin79X2HXoREb3S0kpctcw8muN
7/za7u4LaqXUthhNM2f/XXBpX64YNd7c8hmMortAXomsftaDoD+OL3fmG3Sk3//sp+1tvq/AFXSK
z+E1DyXVhoadJa+Lxyebk/gQXZWA4itqhLbhawq00XCacHAVV5Gve9AsoHemi2zA7yjt5XllkleY
XZszpsLwtHgn4scvS0Yi8LkF+nj5tQnwI4wOAuulSCxxBW+DJvWZL7Nqd65llrwC9jATZKByEWWM
sHXlZj9J/AFPilY7kRp42wRBvgWllK/AXF/Wf4xBWjFf8z8qPnKee+YufSEONPdJUcO2g9Nppcyp
ftxLOb9IBMtKnwzIoBgXZtpdeFTlEF6UmXKXNPjD5XQNy3i71cMxepPT5LLwrX+R5qdQfpKCLwbL
0cln48Hi2GM1lnRqCiHZQ1cw6wM4JLylOTKdtxpkf3O4Vk6JPTsuHnIetIWDyXPp4Z9OP5H9swtr
dJ6ynSlY3S3hm87BWDHizFdTcNsVdOrWXW9tT24JRuSYwPr9NLRE1HokxnFHSq74mtAapnPdUaP+
Qa+i1+LlB4XFN/RdQX6lHaJb4V48j3XqVgLPJxQsbnZQH/wTwXVwf1hA0c+OM5Cni5zIbxnlCgS0
ENuoBnetN3TMLie0rIl2OQN1We3rp6czKxpagVVH7B8s7YUfvhzioLIdVLcYH+Fi31ls0S8D5non
tKSE5CkYuLVgUvqkTefpEJ+nSe3WBOKFdYtQepJ/0uGXZteDPuczyopaFeurkYBkl46FyFHgfN10
nRBZI0f3JQp8rbuxzReNfdvNRXkJvA5ZVM4w+3P9ITup6jea5wVWWwax1VnGp6r5cuAKzwrn0obI
DdekI9V1uUupT2Rj5BMdjtQV6RH8GLZJvByBiMFVd1N2+xHNo04eTgjQGEzADWuXZsFRkjZyJMYq
5sZyyaDl8WBB83DW2bYXBjzc0XKu1iDEVb1FAhMddUuOdOXwqoddLRzydbxWjwRhTiZ4MYiRK/OO
95GvTH+kJf5aNuo1u278/9ZDAqcwHKwrFBCJsrBDzZtbEwY/q+KwHaiUCyQQYS/BhZpL+1sTxp+W
me8ii72t1ja8NUD6iEp8+lKxnwT7qpdC4q52NVYAC7Tz1YPTUFhQeDP6TzC9eEKvqnjFvXD1GS3F
NpJDvZ1GqD56rkx4hysnJwBY6mayr5EqN4oUS7maG4wKr5i8AKPr7NLa/x7uBnKGZeXPKGARx0Qt
ZRoL/9rcAjfOmzUOTIcaGidmqY/fciE93KnI9NVA1aDVkYmeQttoTpDKrySpXVDP2gE9IOvls6x5
jkxIs14isvWCqkRtKEZlww6tDczIhy4aNXJTqFvZF9Aax60Ic3gXfoQ+gYLesiNZWtvR8LvNHJr7
rLjYDqlsSkXuotCFkGqi9j+FpZemogr9Yu0TmbpJ0bTjwzUYEkGZ2gUKludS0jf13ulrq8Uu7DGw
z8lpx5lgh/FimsqOcu0IZnbO1+iTf4HZmsWMSTtX3kV+gta3HyZKnWodIoZTEaWS8ktUbijGH//f
UPsAAIeWieqvO56f3dBx1JkVT/WHuvDy51xbJu4rHsZCbhVbTrgUBxk1FUgAcW3K+dj65ex49GkM
NzavyqtMN7G/YmADRUu6cgYi1VlZ1VgbxSgr0W3pVSr5THix4Ad77x0Q5qJpCk/075UgZJvSQ/zt
/d246YvXz1ipFwDJmb3niTw2U3ajmtOcdbBuFexIDnf+IrrVUM04IYFRrcwMCqmGd/8t/JJMFQbB
KbPBQxcSHpvc8icVPyndlfTQI8dGDJvPEQyiccPLdz4LHfq0dCGSPWrqjtSVeoJBidn238hOwhLa
vDMoBWz07kchTJJLkxvT8Sljx/MxvY6pj8Yxqb0rD/IWfk0IeNVCQtxOUnmuoDMG4TnTosYTt6tJ
mBOPB5Gz9ryCEvHDyuWZsyw6scJ9EK775dQA9bApHNQIHxGXIZakIDFHrXhVSEEWKeX/0EFk7e7n
BWk5NRIaRjwbWS2mZMYVhzwC+5Hbs2MySE0vdS+/dqtOyzlZpVBkLKsYMycPBG9uk7vtM7p42fqR
B6PIf6pOGXyM0HFoALcT1Q71z9E6jCSa9bEYQcQeB23pAlsuvVLSylhYXF4oPZdvEpJ/0UhTWNEI
mfoReKr9rpsBv9hJ3oQDdOxGsXs+WMvF2hl4ZlLXrNuoAAFNvi9/YvmpjwEB5cS8piBbyvHJfEUp
gNfI1hkdyqe1Cw7uScrzpAa7rZ/PB41ybTldd/Ogup/I6CCndi09LQt6wJK3wWy4TNDhWXoko0TS
EmTdLMg+V7rhkqte21LQflj5f1j3rQmI3WCu3pHFkSexX3H6PiS55ESjIQeABBSlSYJBuqRMStjk
D+oY3asSLg08ApiBNmRVc9j9HWmNHjiOzup6VWtjAibp+7WvTkFurgV9jY1MoF0pwb2sd54tiz3C
MsqQUUEsRpRY3NA3mLev8fiSCw3wCtv7eDcCr9lBZKgDo7KzY0ImAST4PHAl61QVD/PAViVA0HF7
ah+5xvpHEaQ8da/ufHBp5moHqFIxSqlh00cAxAY9Fpu73jpKRX2CExDXbTT/dAaY5mXoEysdZ7sB
677I3Li0mMgtvCKgRngjOainxyHK4wjrn3vkjTD/Rzve62OLEZy2NFs9rNP3gS2xfIWSsJYrpWJk
I7GZ//Q+TSRFrpex0F4qDz+wptWbhoCn5cNuMM7CuS3G6yhFlb57wvJFRNdfDMgsSFK9RRL/ULiD
uUaxQo9E1m/hEz96G1S1WH9Rp8DyRQ9+ZDnaD1Ct2OSncgWVwCbUmPXxKAPy73SK6T9Z5fxDR2av
ejCPZIaG+uzB1t+T6Ek24Pky//ydPbzD2dmWRFEpnh3a2l7iKHmh1WVtdsQ4ebwBd43DuGQTQduk
ncTNBt2sMhQWx9mtsrHU9tC8/YfzAAU89RyFfRdctcAqLD7t98ClvZNFXjiKqf4vms44O8NrsJtB
rUjC36efHjfMJa8kGYnDjK7NhGoWv/IKhWg/pC/Ovj2ZGXDAjKOjeA6CgRh7jb+7WQ2h15PyYAer
P1giuWvhLVPs4ISVYuCTst+ckvAnlkyvnaYZEMOPj4/vNLMmvuiu/uWGJB9pYcGAhlgd4vw70Uyb
12qgjMg0xL1HjMJoGxAD+Ztqm6xK21G73XuhD+cbUGFhJBlIi6Ue7HfrOTrVPlr5s4TLfLEynOcQ
P2oGrlQ8G8OE7gAzoF/R1lIfDRotpRivZLVtPx/n8D4xAvBD3F7BMoCCWYQBosDJNS6G3laLuNyD
mFtqRiDD26k8iVjZa5eCElmoROX2UpFHbD3CR4Sre9MCm0lxwd1C74Zb8bJi1/s+6aMiBfNMX2We
goCKgwOo0GquCnAF2HZD+V05/fZRBF9VZhc6vhqLdpEY2giAVGi8hy2J1ZBMkRmjRErL3h8WmckC
EE9LL4ae0nvQN+YJowwesTxz3O8rgcIa8cetkrElZzpTORSWhdf3okCSK7ZBgwZUvbeDwpt3z+r6
9PzxZRnMSvvGL8A3r+l0dTESNOEAFeWumIi2iSsU0gSY7Mz6swzz2P9F8N0YxCaf45Q0MQ6P62lO
JvylfWeQTr7fUceKOT0t+yaVbeAVFHb6powwWEQ5xrNqf0C7qtL8+dmbDjGrR48BATDDj3jWGvLQ
RZZqn48Otxa1rw7l2ewh0izJa0TfTtDQCeWSlQRYY8NYfZ13CQ0xM34BygFMHBKoXtXRSPcqisfn
mcO4ytx0J571/I5yti3F1CJVs9D/6KAvmgRJra/MmmGGVcb05XZEWllnYfILP3DB7w8b9RMa21VX
fHZV/uFtAYBy37Mv6EbiVZgfLHCLyXJUOsaYX2fFW4g1pndGxzfEKpME8pFdD2Znvg/rm7aZwzPD
JsqSm/AhYcF/gv2F0AT1CkiliCyFU0lIYfVCoTjAJfAs9N7twYRRPfPTG4PeZje3Hy8VCWyGf1/g
Qz/w8xPHu3Bw0dd6Y9+3hYqzZt68s23zMCVJYwCw9IZmJTFY7Z7K4KVWZCNR80T9tWFoulKGiPRC
aTccfpILIOp7xwjrJ9WlXlXZabzhN+smvzNjQd6jdxcboYmfrzV3kHknVyXMtc/IrwN7l0eqjOCw
nWpyRTuSl9RoAMpgS3Cb35BMl6mTJXWphEckqDERsAlMZRIbDVTNVcJkN2IWSG2e10ZEA8bZ8AXb
izKLojblRle9o9jUpHpjiHbHZ1TEHMY9soEj6yT+z/jWCQoDbdCUVCCRjfVGfcL15JyKdDzF9qhX
pk8xtNajeYVZgSXAbq/WBMaiw2rcBibRBgj8BbB4mM9A55HkqhVZlBjkHYUaqLz5BRvoH+8TTDGO
EEAx4iQMYPIhrs0xK1cu/VkVEEF2WldYx4hJJ//XNl7g/2rfA9HRKjODpp+f+BbYNXCPXC6H5vQQ
bEGO+Ks9ZFjCRsAUZBjGfZt5eHzte1dOJ8ldp1X/Qy8tQn2iC3QyoY+5cu8rBJMX2cdx0g39NBFL
9OjzTcnAE0FxsWswKEGx6c74ruLeNK1ifEjVmtk/J6CdrZaXy8uczPzd3+5qYyicsV1YqC31adIO
242r56E1okafKhKrKzzEf8K/9SapzVuQHtQkS3UbU1CiadHMd/mWzIxlLTsTyS5dE8hUTgipbQ1o
JRlFw1ExECyTWyM9F2gc3q4iZf60FMaujaE1zK7hDHQRGESZjJqQTs7r5KURokPIKsyZX0hZDEKT
eo0ruN16uPFVaa8eudXFQdnrKeRVEw+rgLqvL6XlaaRYYfxSV12eSmkzh4z8pXSPUXjY8yyV08ve
HtpcQzZtZ1jYR8H5yUSijvDmqlgnW3kgsmiXbtQkdZ9sg2yghmEnFasFSboUn0ecB0IULgeY6GX5
atvIVSCXmA5CkeW+LZ5PHsNHEJOpHEB04mRp/CWahMYM3oRna/q5NXFtoUSXkzb0WqE15ltVTfQS
uUXuOoeC+EZf56Z6nf2U5zN0sRHgBPdHmgUjhkYgS7J340oYsUmXY/DeBaPJDZ+wEEFbkSvNIyO1
0epWpHVxxO2yquECgyGKys39GoHMRXcE2MiW9N6TY097aXyK0nJoLnd6Bi3941NTuja90hnMiEl5
jLFSmehDjwYhQ3y0agpM6aRj8UgDNEe0E1E1JKls/7FkStVC8FZk015KjbRj7A1mcDs15lTU1fv5
aa1Wnb93Pz27ta/+sy+Xp3X5xkK9vS9pf8/pdMpWj5qHaTxlVscTQTZyDQqe8At3nqorelqa2x2y
69FKGBvR2/3WxfWRk7BlDYX+36+9AC1Z9+cPTAYWiyj8VqpyFLZ3cnNmKXncGhTMINKqSYhda2Ml
K7tdUbpiSR2xa9tOlWwAWfoeDnOD/KTVbmlLVUd9t1P/fZGWmB24WDUxpgwtX2lZe/1z8EAexbvH
iz0dJbU3aBGBdBtjAgkOTtlrW3ubXHb8dvoMnmHFrA0XZeqGRBKJzHbpzcRENoOxLn4zlij3oWgt
hbxGwI8/U+MFvCQXDbdWyjBe5WHJulak4Coy2QbU2NUtsDhQdInraQByyefGACqWHCzSk9CZyPaw
dGHEyiHdpdA6/YL9ywjXFquiCGwD0J0hSXtD15OAqaqUE2RGuXgEocCyVSySo4JTlxs6wJc7pOVa
CwHaYRhlV8ctp89jWTGt7vf7aA5jkTHShitOPw4RUWhtIvNEkaecyAHKTLLFxfQoUBWTXqgFMYRX
7eFJRZH0UItT7il0No2F3mvNtbFC1Lp3LyDxbTGfYkbUvq/8qeyEe2Sk9DmgOXfmjBo04ZEsqs67
mKVbDuK+sG+Lq+bKQpzAO5pCxxfr6hq0fsc8uFY94R1OuQ/2gs0hI9l1r3K688Emtl4cRsOXhLj+
UR9g5MS4yYIsB5wmNiNPQu5YIn/Qkjx9Zdr1DxwK1JCUUF5Sp+hX8tjsuCrklMYRajRg8i+aOugS
QjfjGwoxk3wU4gZFtPawLDiIe01egSOlU1aOb/K4E603NvxO97JRnzelQCfiV2KwUhk+xI5/2J7C
Q0re1WWMmXURn3kVS1Jm3tdGP7pQAkepx80ybjBcbX27wdLbFA6UOWrf4c7+wT6zQ23Ladj2e4/Z
oMI4BN2rWe+dh5CKYXLtxK4OvaT+fFo5FV1mM7LSBQ/67z263jGfdJPNAGZGHUwHJXDOQzd1W6il
hlMGDxnidOBooB+6I1fwPiCpEC97GsK/zbqjeD11o/9lHr/vhsogaMkG6tPDiYBjXV4pzgZ1Vbr5
vIQP0ac16jG/EEU/BRXgm9YzRITp6UTlM3kU12KsNvDqr1ghlDFi00ehFva82BG3ofeSydQIXQWR
/Xin+uZI2NEa6ZC3IDf6CYH/C+Wgm7BmomMKBsTAA/ZmzvtB2Q97gGNTfX1Le9pmq4VoS7sBN+dx
JQ85KfmVPTct88pAsR4lYL7iQCTAzEN9Wiws/PJ+n/FIWxmQjkxY/ArHBer+FITKwYiX234IQZxj
4W0VgVbcSXXJo7AfVkoAIyyBey7ZGO5Ux9HtvA0mSHfmyM+J3PhMA6WbCgHJrumbWRcWE5dj7zGS
4xMiY/EyKYrUhkXs9uniRCfTDT+XMfe0LMUsXGyDOrQnl3MQ4uZxNX0rXlYZ0EOToLq8EBPoRMhJ
HsVlfDBgRMATZfdtu2Now78O1UeMV1TqgfKmF5g3LSjZl0wMInlcslDD09xgJXbMmIY7xGNGvrm0
fd86lM9Q8j1MGme5yqth9qfVDTdfXjJKt2hJv5afHgAjL9IHZeSZ8FjwrH/+vFK/+AuBmFfQICcQ
FnZaUxhO09YPHhdj4rNzkUV+0WnPyfRZ4c51W0s0KKdeb9lxma6BeuKYex/OGk7U3g44mFRmu8J5
7QACaD740E/Bc6JLJSKW0nFrldarIQCXufl0AvlnvrFAwcfBTStWwyInP8SXmqbWvzAv7nX8ACVo
9nzUzWLY2ZbXNyiXhJDOfSyLuwU5FqUl5/eDH8ZGlmYi0Gz2zyj1ou+qYazw6WklOx+Gn5d7SorX
vmQLcC1fC2axVCL2tYhw6YTRPkrAff26iqG4Zr814F0JBmHvEbCEfxJAYA/rtbuNPHl/xDxoP7kE
dDWdRo5+QTjtTLQjltP87z7tdhrni0PlMPk6toiv2bnXUmQn5Z7L/1wp+DFDhhx8P2JKY4wessE4
syrePKDvZANlxmRoopWmCK71xj9w/owFSZ2XiBlo9QlbNXPYG+ZsEQBX2LBaeUADC+GA2v4Mv+j5
qP6hcq3lN/RcRMIjg2msAQzIF/HQdi6gngVTrUJKoIM6/2PTrrTe4cOsohYJU/fU9rXuOPdZdG+2
QVxi7OGBMdV9qa7jbyLHtQ9aSNkQp5k+hZNc8mc4OLNxfq9r7FC6cY0SnkNcn1sBsrmt28CmASGW
weqCVnYR8w2bafi+207G0wafDpLld1o63xHYM2X1xA7UTzY70aaRZkqpc4b4jMaJKGPzQVzyRuaW
xvpphwBy7E+dPBzfx+f7ZKwrweM566+wICSUz98+LBaDcovHjb9vK8ZvFh42MswMY2OXGZH6OBFZ
GGcPKye9yRM+bBmXfIMS8wX2W8ZDAxvTdnJumncv32lPcYSzh4q4e7aMlo46AAcExe0kjnnL/IT2
3h1S7TL1/XBSrteGu+ODXOn1FEQFkNA0MMECUFNm+dAcn+pNisZJ2w51sB6QRVc++uowr222LqBt
9qo5NtFHiDGu5lxt7Qz3HytUCfdMWXk7cKZ7RhKnnGfV6LzQnou0NOTDyPouJJRM0KhHFEmhL62l
+KB5wdQGSTBG7QE/0nmAXF1Fu0yofK0J0DBqSQ1q2nkns7CnDtCJNHuM8B63jv4Sj4eIqkoCnXpr
9qAZgWDlNJ5dsbB3/zVd6ics/0He0ApK09Cmg6hITkPFaCrjJkehh5ov4LOrQmoMF616HNXFynC4
OPbZZNeTDw5BUCPr2Hbr16RPR709Hal++Ywj/GUOrlX5lqwAM/668HBuPgdVMQp0cx4o/B9haF0G
F8OL29L28DGa3sqHtCIQs3l8QPGk5fF+wbzg7TYeC5PpUa7ljqORD2mbommTn+t2GJP6mBIaahfZ
+ftozhqv8frhZu9XhVQgdzdtTB0enrX6dt1tuGGKc0YlWSg65/QtSl/2CdQjCCRW4Og9XaclidcB
8V9FBtnRL498d8pJtJZpBqcfmNaJE0SQ/2yBXUHNY5vwOnhMGoAheStQfnD93efE4zF+Iv+XFAKy
yTXFmHrO9rWZSktGU4YzFDgpmIUgfkGVeV+C39fBrq14CyNdexJXZ5Nv/DqoWDrxOjmKY/HpWVdC
gs+EGatgTNU7aSnLZGgW7BKRhO0kjmdoPwMyHLVDjhR4hK4wFqG4cPikMVJbRVZc8rJ34ZfXQ705
LsnWl2y2Wd061VHgi7d7sHv6Ki+Wvi0EU1iHODupfiqdIgj3PbPnVQOud08dt4AENO+dIBmptmUn
DvO8TNpQABt1DsG2e1/VE/aEktVZGpFhtWlCeMf8D8MMu5IeEpUddkXttWSCg/pFqdDH5wpdSEDJ
LUSauhGeertfLSfTNre5cJAnJxcA00NlFvjco7/B7Dv1hmMHaKdbKIoRkz+IJbWQ27cumo4p4qoC
QjOM5FATQ+s/BNx6hbpQc0hB1jwxtQY7gSh5ChU+RW0Y9+hAzwU/MSuUa6tnqHHnOQes5fPuW0rw
aU3occ36FSZflkbKNf2hnXF2O5xgdbgNqrd8Sgd5aJCQQBnHa2CM6qPHkDN8jZzueJzyrgdZvGt2
PiZcfRW/WIF0RVymElHiFztVh+3lksVZ2hKfigrKZSx2O16QuSXMEHz7KKuzludLew/Zp2hrtmjv
+BtttmFYWzVJHBTJvoutKls2CPlGJqpeT7vIx03Gp0lFE4R8cWg4Sv3CdVBnBGoukhsXROkI4yOB
dpMiyXBE7ULcX7p9nXmHkCrGxBgXY2uAqhZQfFgG0bs0qhUQPL76LxAyTTnMRpIuL+v3l/CpVS7H
oiw2u5AKDFh4IgKI0QCbvCeZBFT4/nWa3rlSDeHYghFW67zaAjuaoTG6VaSjDFvj9A27YRgNZvBn
MwD7cmomidFB59ovZK5wj4ghaZPngT0gwn2qPvN9Mb9w+F2jbAGftNO4Kc/yBgWTITOVmB+zA48X
d8NJeer88SjUSq+NjwRynDawr69vLTUBQQWo3l/iZ1hndU0oqS7/Z3qisIIzN+RXqWQ+5xJuDnon
3AQ3HVrKZXGuNIbHtOefnWoqeJpKfcj6SqtrjKNa4RuYJdKfLgK6W/uuxfn5jkOo3lwn6yZd/wJA
kYaAYCCp2VjGrgGvtmwUEGxQ6BVfphcra1N4JhQjdAZCjFu7TzgtPPUFZw0UUZBrIg1FLkj762wu
k2TifMGPC8DnVdMmbr4njR13Pm6Q4pcZ8/bitcb/9TMV/smqrQxXsaXKhXPBYO5E7hA01RqTJ/EI
a41Ngx6PPDALL3Ldm5EN543CD6MB2duF+sW8g7wIVKrr+jQGJvYK5f3KenW7iG20K/M/UelsOhtB
bzYpPGq5NcbDt50DruXfMYl10V3+HWwQ4HCYX+SZgBBfZ70L74Crr80ERW6NdS+JcW6Jkl1pSgP1
jIe2/XWypFddfdkNxXKjAXePUcVJaR/DZlP/vg0TR2lm/udqJleemQjT5T3lnxWlpfMhwb1OUfvP
F4E55CK4n6kuoJSvdRn54w3d49XSB2yQcpW80JvpG1LoG9ISNfr4Hum/llZIixhNNAyUPQL1OQ2l
l3DWXe1nHjc+NiT4IhoQ4abMdn3RKbUJU1QkstgZXeZIFu1eCDflfBCBxX645PmBCo9xcrkuZiRz
8GC3gtjt7OaQAT4Ho9gtYqGgSCabuuCCTdgy1XFcTulEP0vTHZoedg0Bp8xuNswtKq94ad9gavVG
FdvqCbAA84g8cqH1q6zOTfc4R177khcO0xP1928c5gvg4X0eEm/O5mZfntxCvWsjKGk7T5Wv81qE
bn81qtaUX9G8SbrFMTLCAmek+Hu7S+PUKIIDCES5tkpajIX3JJOwbrzqA+Ixv54LqHQcOrn6ghBn
LU8wXGDdj57cxLh/0ot71pJ1iRH2H4+UcddM1X303oUspurYUT2cEdxvCFXMFqcDC1hWd3YlwQV2
Gmz4OZFS9UYUCBFeRM5/uR+cvyukchjt0p0XYK1Aw2whDxJaNputEMbfmjnPnNuZJH4wAbjXPbLp
r5kVOPuULp3axqNCdD6L3uM4vjVmd+QSSwm2xS4dVdWB+YYUHKyi1aFASBQdnNr90f80xkF7TX2+
lO9WbxdQO3lSxDVbsqSItqEEGTKuQSTBrpe/ZTcb240rLGdC/n5y3OAQBsjy0ZxebMpD3d/prQLC
LufpeL2aZRLXm7nqa6clD+ptG0y1FANYNzMGZrcFagCMIEYHMx4c7bVz8hlUzRcgBDwAFgPlWHVv
SmhAcXjxoqWH28SRFeMRrKqk0LvCfshvZuSAcCVZJ7Zr/385QySIrehD0ikINsWYKT7PCameoB1Y
MGtLZ+fa0FW8nzLoSbbzgyX2qR9kXTNqz1oq/Qz6ViDDn3L3HqEJq8lGomq7mJSsXy0mWydEmn64
6DALKY0Z+6CepJ7CnW0iHja5fxB77Sp2SyX/DXZmjQa3mr1sgt1sMAtRDBIr0DrBNs9C4wtHsvj7
5yVmcMU4/G1XFP33INTz9PyrE0LLHaFsx2v8U+cPObCUfMC7VBgxOm4a2XcXrUBLPon0EE4JxhPf
D+0ihr0DNbqrQgz3qVayxl/atDwXgA7QlXCdEf2qY0HMRJYA6bZxIdoEj5cvuGC/3r+piwrddUpQ
2unDyvN9iwpGBo4lYyvOi5ccGgAF4bhNKnhqxOFrqHJBOmmwJLDCgXwUrRdr0ZndDyQj3edZ1ExR
vkJX/qPczlzM8aZLoRZd4R6FdaHcf/3k8raVLfw0Esb/blJ8w5tGGlaAusjN9Sr90WYFjd/9rgBW
LaqgsGdedYFShOTHjaiXENUMBgkCR08iU6ijX4RAefE+31nXFeOwb4EM9sJdjUgp8ZG/BYdS16Iw
+tJWl7f2qnOM45yioHcAHBhpe6Bx5QGhkEzL6145SGEC0xArwG5CFJxb1rHCtHEJtqaIx4SYv4Jt
TIh91QXiMQTFcxSqdRY9H+qD+2zX8RycEn8ulYgvezu+mpAiqdygkQf1peSyMQZ1t73umaAsDlJl
hdGIdY3iH2jVstdaVkQ/S9TbE5mRQi3BLU7yYmA92DVse8fvtQw27vUrIF5MCy2t5YpV97owCc0i
h/y6fw68Z10nqtkFlHcZ93bkTkdx3a5pdlbecZJ8MibJgqRkES8BrDDpDBKxAQSPlcZu73hsOOYP
uQG/RjKJJw3J3WJCDSetBwy3Ki2o7tqBqphiTT05PgMAJH0r2ZtzX+ebYy3NlV+XnQUhLidPqEd3
kG2XrTjPEcSC6CLiynJ0pOTW0XTpKPkVCxDhd6BquzPlgUyv8vspktf8ZhAD/3CCZlHQdcyB93d8
Vofr1tQ1a10VNU0b/Ur1hXGFLvvpJUrNAka4VcAW9egDvr9mDgkxisqhOnkXMhHJQRtB6WNVoJgm
vWf5ScZB24xeTwoEFMCrs7OGTBO7ZqdQvX8r9IIzf5nqGsYDd6iNIhSxic1AvG5DLljaBQDNJBYH
SslLdRjWuamTOGeXs57Tj4mwAqMpRjWuGK7NlqwcNEtKhH17rdNODoo2tmpG7U5+IztaynC2AmTF
97KcmufY5hQChP5DeIq9SqOo1KXvhs2bVvyFWrBI/dxszPBLnpleMCp63bPu95hU0bIBAw4gD1Gx
z+4Khu70Kt+bqIZ0bs2gGvtYsvRrVyFWzPYAPlRru4XUE+HMBVGOrt2QxdC2h+VGThZBq4zQ+2Fs
Ol6rsuYU9718KYgrmMOPCO1xIyjKkEbOxkTr0Sx9FBzgbmkO837l8uZdlnHL/DYViAOkN6eWvjdw
r8+WfetR6Y9rD0aoSLbIng7LNksgSm//58l97Je9VwA6njO+fD/JjExGMAIpWXW4MDkhimHc7yD0
xzgArEGSqs7j00XONIAyEA1+Ypx31nhkMnecmeXuztURNmBT5PWoqCkyPs9PszcC8G3JNmvjR0mJ
vl4GGEJkdplCzgX6O96OET4MT82JRomsikKh0g8exLMkka/o4Ky5Xy7ooTdD9tzSc5Fv+cAuS4mK
0i1gt5N7cKY5Q01ox8oMSMOR4Ar6Q7OaafTAPeQX/Yij0UwPw8TsPeDY6Ij9LdwwCxqarniqpJXT
nOGJFWOXuL3HmU/2Sc48vaF5gFBOI3EgBlS6SuSxI0fnXPUAEKTfQZreLW/gfIbfEK85zwrhmriR
5Q0eCwoRO2/qS66vef6NgeZMTwK55xzDufp/nhKmwoNgb49Bd30DQtUitLj6ZhUtoKGERoK19gcD
mgIS0kNel3vMWWGqVXbfm8Pt/vSDO7+C7ZigQvHWDHuxZ9ftUgViSLDwNAggdsy8SsUwE4N0aXdf
NroTV2RcjPMvd9mU919B5n4xCb39J4LHRQ5prGAigJI9xZfZOos+JoQmcMxVAChg3cvlE53Op6Rt
hb6m69CGddMi8VRy2oI2bZso1twskix1aB5vh2GmYOvN+qrTaCvCmPJbtithFlFyqdVG2AaL2/Mq
gPtuUV33to4eHok6zbZxq3RujxyicRyORMgqdpv4rDLs/WJJCu+R1WRe+iRlXb65/2vriDrWCZre
o+dtIdr/Ep6weVAdzqOUJNM/8eUqxztcyt2XPLMIvudEMkBgLaFT7jgNz0LBgroowmdWjvsIH5lC
9vpOfDNfGA+c4VlZoqnHlthBrVODuArUkLt0Y4bcyArA/IuHpReJwA/y3f5Vbl2ZgCy+roZPUD0b
m78+qGk62P73Qaj+Ryp9FaHFZpDbwR9o4jOTCP/Jtlj/MFeh9u1bXJWK62Oj4wtv/GheS+v9uqqr
aW+purUjTANZDTENqVFYJr+t//1znkU+kLFyR0U4Fh/B2ofNbYMdpXT9BlXmzFw1vaYPvutx1YIJ
kXRXe59hek19iwoA03P3RGKUQMwObkRLs2K2BVH3K8F1sxacQb57F25EQsY7V5GIA+2lXyT2wI5m
MOx++ooFtxuemLcFvAIPAXbDtDzfWM9EpfHwkIMhs9h9IDoZm5v7ScnwIXeY6xAVdo/w1mM++ybP
pBmzjcIgSHx6wojaZvEsrnpfNkgfRzEeI0Cidev8x4ojtNPCqo+YcM6jWW5aX217lpVTn8193h0x
3FW+3UGXtA+Kkf6WPtRgkOuyhz7gIQeFpTR1i67Um2uY9KvCjgJW5NgssvNAsYqxzUWoip3esi/+
EZ+E2LsB1t0/6pWRhu0h1DRpljadEB62TQY3h8iCsWScYHhHcJmxD17CwgU8nASNHsrKarYvqz57
TyjJ6aBDD0/hDMR5aiL2u15Q2u0FL3fjUmnLV7m5q7QHtT7AUjAbhqSulU2gSYHfyQKcOosML0gk
92yuDaABtGRr/T5sDxrbFfVomY8wqCd/UsAb7MXv7pplXDIwaKWelP7NiaT2lwdt5f7s2hGmIDyd
4aFxsSPKGp8RZ0H2g0seWMxTrgFkOalpMc8eHiHWxH6sWUlcFBaDPysqeeTWxKWtZU9ZGU+r1pq9
/3soa7M1Bq9l1eqKbFZogBKORu/dGJu2kyHJfXRZyC4V0WBqp8hq/9uPYGUI9PW8J38OLguDA/o9
clde6HY+fJJxC20QcoxtgvVixS4snIVxbRTMdp2fCgFJK4ve1bM9tBPi9Eq4P1z2kN6ctqBIGZCO
1h5erw7JCzr0VHELMxKONB3ifRjrLlf4j0/nRbQlLTDbcWDUg/i0F2VUKV7fsnDCa9lhBm3nu8Nh
m/Sv+VrXSwHXos8B7OmaD+y9JJwc5KP98oDff7cizW1BaWTBKsb1dQD2PBFK83T0pLk41dMOIi4Z
+zbBIQyReHgze49xgM1x+YZZubeITotP7xfDDPQR3oZMY5VsvP+5P4aZIjoWAqbuELJyeEqS0Zwf
8bK9nkz8CdugC8xdnpmRdkogOGsusssRrnf8esxgEHZr4eUcq+N7EoMzELDDr7Fceg8T4+QpyLA3
WaS1+ngkPQxs/FZU3wd97pS+fFwkEpX1eYc+zk3vx0jDmuhS7pvnew9w4LGUMEBY3MnQQknIEbDN
Zx6hM1O+WiuxPePPNHwJHhtbD5sARYs4J8WHIfQlQaAQ+gLAXerCTnFpHEnDtOMY9gxyIHp4+iiF
Qbxvup4jiWnCG4HrwzhFBb73Kg/IMdbMoL+gSN1AapoYwra5MSGZ6Ua4cFgTlzlxjFbpCGXXXCBp
kbBYjbJveQgSv/bbsN5YHT159xEoUt56EvHWHEexnnOVS9z4vtFyDCz796cclPEkUQlLu6wo9A7K
C+ZUM2SotRZADAYeuC1F8SNb4uJ9aW01n8uEADZRq8fBGqNSu9D0vHq3p6ULdQTzaCvODXtMKTem
WAJxgy0aQcbBwKaUL9pvjx8p4mGdR6lvcTel/nmAmP9a63waQynw6RwF6BZUubyg3Yu6LtQDZiTg
RPQ2ovYZfn3E8TXKRhhB2v7BkrB6b6Oy6C0P8pK3zfumqXH7XtaP7TdcTAOYH7mvCDqtIUgyOGoD
AiyPdCZXabfUtyTG9Se12zuKlEQE9a1hHrsxTTW+HxlVjXj3E+xnvgThaWOY5AGBfCuhwYk+dfCF
K939BX7bJdBDZZY38YPKLWarfbAlku1goW0iiKO6COLCEgi5T0soVb3KEyC2tG4M+BQb0SSRIfZD
tASi8QpRqDcKDnozbPgzo0P2/7F7mde5eE37dVDyrur1nd41DLcmHLPJ1JNqMHhSISfLRaLsEfaI
c8NDjb9lVOgw/lkm5He418m8IeVbX/JJYqhBrBbDNljGGzvXqwf63Ej6lwFBUY/0HZ7TNIBoqdLx
rDizMrmf0jcQhXxW39ro/NqG+izO8UMp30px7oZHSsLOpZiSiHe06KULeZBKZXSXinRM9kn6aJ11
Z7I/dDsKZ217+Fh0fLgpoxHVmDBKlhc6N54krWgsqsGh3Kfjm71bDdTFFI16D6FZ1fHUvJTK/ajg
AjoNHzqHGi72yDMa5F6QTI6cVep2oVCePcMp7cWEegNlXqYd+86SongM6N71B8WdUcReKsnklRLn
1jFc4ZszI5s2gEgbJ7xjD89oM3Vncu4hYcDTm7i4NnlMOGCmDnfan/o2z+cnLKYf+VpjGgShCn0x
96Z8Vj2Yq4o9qxJpzzAbW46/RNuyE3g3pYeC9HGfP0OVUKphnKEu220dPw6U57khI1HX5NTXJzrR
g/ouvoLBrjtv8eCNQFuBo5MFNVTOh8rI1BX7x7OQnaUtXb3bMnp2Qve2VSS9ZckwGqndrbiQK4AP
GXPuYfv0CJ4TZzMpgd0sGiBKVJaMxxtN4Ll1ta/T8ptuR0E3ZYgYGvYpAXxn7qJti5BACCzf5zj5
5AWUWquNxAmaGhyLULXpZ2G/6paI4zslrlA4YvS/b9g4wxhl4R7dZZDlS1JpxWx7UKQGJuzHzj68
x7s89bcTHTHywvtIcB8SLN+GgCfyyWjAHah8lv1qvPRiSkQdI1TBXZvDmRuwsuZaWuTrCjbRk/qb
zIv9VI3mgK72gRrgrAjHDjuiHJQ4+qmFsdYNZ941ismcabP6tuiczg3zWvKThSyWQvXv0Cv27HZh
HJ9xbFbuHkQss+20CltZgtMDmGWAHS72MtJ1yFp7xnxgV/EyRlkAdL0qDgeUN4n6SXJs4UoD9Ywf
VodHd+UZUsWfrzGDYrmp6FDIDmIIJAWoUNx+a2xBT9SiHO8GGE1e3KxmcFGV5cnoOPOVLi8ZKA0E
WiY52yWletZc2GLS5B1X4eCnjE7r20LVo7kpg/pv6WY9Uh3fja5ur/aAnThZcizpkYRS1HP2MID6
+tzpUsxChdAdIpq/S0h1VtkCizP04QG899SwY+VEn8fyxbGK16MBSCJy2UFfv1Kzs8at0UlnxgeE
SmcYGjt5mc7hBlh0XNMn0qO+DqEv5WpaIcs5dajCfnisDs0Zu6BHHnvsEANjDMlLMuyAvh2x6IZc
r2k5thrhsD21nrvRIIoir9YQxLAB3pXzCzH/YCEbfp9LpXV182m3wdxmIMdMzL9A+qvSNIF4FRZC
7SqTpqan+lvdNA8HS65FMacyvAHUH+r/7CjGOawwBgMcz6UEQjwW4DmF1IVrfkMass02XMbQqCvC
ZE8aGS3WIiAChUYE8UKmt4DWUJB85KFdDzX1i91FBqDS3lo/80AghKt/66aRmVxKu/qlhPVB/VCo
tK8d+X3aKHCGg9spYqsf0Uk5LJoKBCmOFliC7ZZG6Umaf5JTEAuPANm42m0r5WCwL89Tfk4UwQ3r
1uGqs6WkMvk38h7VQFY/jaCwZDn8T8M/O3IxYa9FKWx+8Cmky2cNV2BYb64gZAkDno2P+IKj5lMH
FRGJWCAVNgUwypVPgTlClta5Kj7nKnlsbFr3R6ricP35BlyUzv7++6ZlDm46/Req7y2m+C8yVjTO
xPuUwqANzI/HiU1+t90/bF7SESzKZDQzDG7FwIEgBNDMn4QeIKf7/4hSYWEqwkiUhp5Ibu/Ez6nq
XBHtqeFXdeMdIfX9syvxAk0mjWeNaAXh0EvGSk9wsuuDtQoxdzt4GFGwC5+Bk0V7Y6vfLGUxhrFx
tlhkyn3gE4oxzB5Y047dmAQd85GCjzaY8jAwL7PN16BQwT5+fXYTqC4WNtVT1CWMTdqpTR4lCcL8
467Mo8LmSOBkjfUOGlaMR2Q/ebz/4gxOxVfQd8b16rhG3tr3H5X2i1Xj/AslH4JBIDentrKamvM7
Sqc83eZ6rRAVNOuZNARxU4l2KPvg4TmGT2cev/73c3LpmBg6hv5Cn606HiNyPtFWijbuB2CMQ3tu
YmtsFl9grJM86AMyCLg/x3TBpmL0xYXL2zZuXpTAMsJxk3f2YBo5DFCRNLYv0iFXDm/QAGGpUy97
sxfdwDQ/NN0dS2vI728kky9jk7K289xq/7wEUCEFkftpOHa2ck/U5E1XXPMidFeUP/66AZEJZfrJ
pXoCPTR413cgnADC8LEL7d5L0OcUdsZfPjfNmTVivvtFVavgkLZA9L40UfeP8ZT8rWu7xMNnokvj
97+5KR2KS82fjg83ROUpgNdzAWDZmv/Om4rY8AJx8PBMnA9m2HKOrYekJrtNRhbra58KwvxTvoqz
wUUNSxYkoovVnFTo8qjpdPWkNBA7is8jaQebsu2SduEDhaq68zf7p1O1nY5d/MlBOXkjBY/VQpXB
JOm9baTl1QhpLAL3r1892OaV5XgkAAfSLcMZMiP0Mq9ZT5/MSZeOuegpA9x/mvxb2EsQaDLBFGVj
H9T39RJZ7Kw0xN3EELll9rcBQqv7rRE9NEfLgB9Ez610TbWlsDVnCaiUqDWlyZ0DQlsYH9QbkTn4
lEbk79KLBWBWMSVXhNrXvsVzeESFQcn6QipcasPGqPOXk8i+9DxGS4AS+SKTIfD0Xf8b6TQ1JNk6
DQohQnr3xUmzgmQ2eVkA6/cmHnyRU9KwMdQVxWP/uy0CCKY5eLxaDdDyBFBTQDLsXRDULVakAU+z
+j+XtpYUXMGPtKYF9D05jS0DpnsLJj5Cic5AmSbvJWfW9Ncx0b70XEZG06Fdnn2Cl4TdzknukoEe
MLVzxTNrJeAChgyMaRAOlBPZ8o5J22uCI+zz+M2EwjNepVwAroKqCFprWKMp1DBQ18a1h0CJrxMP
TiU5JOo5I51yMuqWOCFOCyvLUlTWvVA3vg05IbLWDUzb8/qK0j23i0eWnLER93khtVWQyhJ7rYpl
JZgQMcFN1dkEvnd8UnnWvOx1mq0+EITgfuUx25OX6Xrwne+6lVFS2ZANvcnX2tOs4WtVlGv4zBpu
tzohdoog0rPc2JPzoEwHWHR5GWtI/VFnZlCjL+EG2Pgf4Sicgr/4xqEuH0v71Ti/qHMQdoePRMYv
oUN++kwndpLzBkLQfbc/7C2L9etIi67J9h16Kn8QlSnF0t/GUHTh5D5qQM3wgfNBcuyko+/Ivjka
mNH4KSM8c8posi6twz3bNEnbJ7ettUZagPDDF4VNF7/x/Ls9tRekxmeXCZWm51Cv4Lwpmfl8U7tJ
kKetPyFqmXe2Kys93rqUQZPdRJyUj1XTG4sy0/jYZ7CjRIq3Q+yZ3aj4i0MqE3OtQpa+WwdIcd0l
GiHS0pZem9UDZOcCKgR6Hdri6qooiyLdZUJTZDf9HIX7Zr3mLJuAS3BOxYmDsxrQDsXXrReEWHp3
gMlhp2D4MMruXMx0Xcg5kzSb+2CNppyMWokQ3qP0SnGSmfkQVS3nMrgYROeXe5w1fadcDMcfP2p5
ycVigDwysj+YMXleSNTyvF9eEobnmZi9gEjCSrwYL03IAE3AXj7zzvynb1/qS+6RIH9yZfqxKkgb
02yA/3pr/EeDtcv0T9ulMsT9i90jEgWHwzVFNbD37A05EsAGO0juQjIAILe1C9W5H2cdPDmK8hbL
kfuxKLlkI//R9yT++MiwRLaI6nnvp2rI5L+LSQWdvGiY+mqbB3aZvU21CnmUMvnRBohnT5gcTLfU
wJJEpJknGWXDtiASOcLZNE+EwYi3KPKJrFfFUoTodUwRmRblQ0tybxGPqSTwbRBVbf3n/qbJpdUL
UgibAQtSBGVOMr62FD+mKTsw/wa68FSmMHX8Q5MFZkITaXlk+NrpctbpmkoSg/5h31qB9w7qeCxZ
ot7WajUo2VeBypuqmNvv+MkRqdHu1GgHGJZQkARaQ3V0pvXSsnKi54+NwyrsVMfuJzfKOMBins4V
z1E6EdGFsLctCL1vj4tG6FYLxMM1izCIe5XfLYtRHz3F6fmFTiflHyrYummLhdJxzANEOLVpgXMu
QCtnVkUDuB577Umvrd0DPCGL3WadtjOfAT5CDvG+4DW81j7bDZH0OwVUOx4O3zFaws7yn1LrF42i
E1AEMGGqUJMfo0Dt3lkj/X15hSrMHYisOlhpsuA/R/QZpSbCXnfov7P1TzV5oKiqC79AP9MC9rru
dIlmChGDG/ELwyXe6HQwOgTXhl9EdB1p0dnqmIsYeLw9PHZHW/joSVxx8oKtVhmdBiQ9DOHV/Gze
6uj/EMd9bnM36pjzxBuTYvxA8npBX7yW6QXkgHglPJ5SF3hmssXssBGSsTp/OJ3DtabpPENKNrhI
3u20T77v8MNG/5qDH1dT1++j84Gmv9OZvwDfOZqw3WnUyW3b40goY/nGuMW6auFEFtUZWobIXZna
sdNIF6V/4V+FE/4dvEkxUtMQp3tyhaEjx+he+QGo6Xayw8ypek+9y74Ig1k7tHr3X61mOD+utEAv
bsVOzYR+s7QqOIqhqo3uZflVb7gzhP8Ng6H1nNM9UKRw6ScbAttbIvUZNPGtjKKAyGXZ83E6kvkb
0JGuspe9fPkDXVYLmbVAqyfoLwxtxtDypurhLxoq7P8sh7kPnlzAYxhbz0yrJwN81hwKgsstlO1i
sYBJBWOb6oaVotby5dOqShfxEny8NF1z+w78X9ttB7kuatt7KDHtEvezXb16rcieBV0ZC3u/y7m0
v6S7FRIuurN3PlK/jfb3VKF4gBm5uQXGDFmayW4RWajK8DX3+9dVFGh+3h87HSeVzkcH2n5825Ye
x4MBLgocePt9gcwcoz0ISStEQ+nZ2Ryd3lI1bEQAxjYIZSSQpovPIt3DuBo/Wb7rSEgXVUL6hVIe
BeRBJkQ68u0FyuARFzzg4zxS28hAoZUvf1Ho1iZL84B4mPQ2Fcj6DMmCUFEGOePVxPfn1I7mHsUy
pOADLp2hNW5FmMcIumK8bhC6SVL8M1vgbSNGwEYarB50b6n38EKhvsKNWzLQOiuKwhChy0sRp9op
JtUP4tMAFFRJ7f9SncNrN+DP0aZMYNQH7L1JvdWs7R+clsX0YF3Z+723twli4x4u0OHo97B96FTd
ih/ltFU+xkmC96RnFINnBHGAHa87fWVv35GyVIzwZ9zshW56cNBPx7XyVMwdu+4PQwb77y46snQL
6zDcpfMatgHcQ5kBzw4/anvM7S/TOuifSg3NyZE+q6T4nvUeRnnOP0fHQahgUXHJ2qekUrnY5l/o
Hlr8uuCFTxwXUrys/kzHHAP36b7qcQn4ejG3bm0q93GHpAoEt16cUo3+LoJQG/TBpcoPncWPQQ0J
jrvcHN52IX7u/96J578Fg1mhWr5HF9kqbOr+fOfvQuH7wIxqLSGmgwY9ork2KVhAmCfZKI5Kz3Uk
1Lcw0Cm4o90GSi9KGU9povBKHB9z+WOaFW8xmd9zaFF/LaagauHx3wJq5LuPCYuPsK7u1PbrfbmD
uhoGLETD/1mf8Zde6DlZ26cR4wy3iV/2zWAGJbIvT6nHthb5U2DRP8KxJESyQSpBr0IFobOH40fz
CIzkgBzc1RNFKp3EDqN9lWtC7LtF2ayDGkH544vM0nnGc7DHC8L2KQ0MjaSy5pgcQRouPpew1V8A
MgraZwhLIyJJ/dZJUfs4zo2z+DwTrkze6zfgKc5DhTNRjCHYl39yhteXYxKZhtt3Zs7b4PRlpGVk
VXvy7lbFl/VI59k5fmdChJzpII/52Avo/Ln90rJNLoq9DKdHrtdVBBvSsr8PhQ9NmsgkeHgy6uR0
XpTYR+8OtE9W4sgW/NUoDQcs3izdoi/oDtfo9DPcM+84qFruhUIT2ThjguDTS/IJsmrPMzLe5VgP
d9Srw/Nm5XGcG/wkoRnodgV9MKej1PMk9TPaMxSoZl4G84hkq/C9XGdzgMDjimCF1bmUao7M2LWW
DxDc0T/okREIwoqFnhS1u6EISlTpUa/RjvFC1olgfmJ1Dn2sSzt4PywFta6rGICgKqo+LjBd84u8
x/V7WZIQy9IDntGeAISS1x0dbwSmJ/bT8pFapEkFGqex0Ououh0lRWYvzqvuPYf3C9hD3X2bowxo
WQoAV2xDFqrLa+a3zcYSGoF4GlwOVQ6WoVUDzXdMPa8tRT7lFzofGjDZuEC6aXpCkEkxZc8J92T5
ak99GG4RO0zmc8Sd0H/8efP1ElKDoq8SSzWBvzrzkCth9iB0UcXOXKL9U7V+DPNp7f75Js20IkAY
CANmb1YPvqlOergHaUkwePvIIzpiLNRtEDrRZEhOryob3up1kQQlmhbvlY/URLK3NZlSi5JACFuW
uYMIyEXWLQVfnApJCXbZ1mIzHXJv3oQrybPkWFc2ub782YB+fc1lWkQSMZR008mByMQ534+Y7cOD
i5LEas7OnvYDTKtOUFO0mILc3/sDTZbNMaUmt52c3OvmIVHeXvOiVHnZ9p4y9bcnVUeePPDcVgK4
vQm4PRceIstzSePObRmWBZ2mMRpR7UjrKsS7ub8IpWPo3Huauw+MiCt8f5fP5Ls4aXLlWpM3zza9
j7RLM8HB4l07WDlruGPsCEFiMNBM7UR/iyKOvc5ujd0UioAyEjWHlrGZAex9t5TLLL0OY//BmmO9
hO6s52YLxLWCK236z7c5VtI1+qj33jh4KqnRf5YXXUu9fS+vOxXFf5e5PvAZTtILwd9tPHZ2Lihb
wXIIbLacJ8GJgP2BTPw9IJWaNxWhpc4DTnUc9cTfHEXOSwKeBv2GhEZTyDnu5AoxMu4O41K7OCHW
sVPOLp3jzfDIO5G5MLRheVQrRv6yk7mnYeoOpg0PjJrZwIBZOBR7z++FmF8RKTJq8nJzhvWTjk4f
brQ3gT4ksF0hZ1Lsw+oSpMt/5FWh6d0AXVvZ41KjO73aCKKECcyPzn5dSZj5wPnOjSPycjkWHxKc
4sFl8SkBDljs/CB8tnbTjkHZhsA8JO+F2SXyGCtI/uSyoNdR1cF1hpPPs9KkGBavEq2wGm+cvRkx
9AgTanXD6sd3OPmmq4ZKGXWXXyxqJnc9O2V+wZX9Vn8J9EocF5vWdaO2KWPyCXGhbQv3t6EvfIja
2N41kbvQqcIDhKp9wYUrLMnhiE2sQLlDmkVYSx/yFA7bTBQTKL5f+5yIWz3mabqrIPPohY/78dti
DZOQL8giCzJVd/0AwECQ877aLoG+SdUFqgmY5JoQtOXANwVWo+jIDSF+8ck1VetlJWDtl7UeK7jg
EG//h+QHEPW1YJ1gzBtopOcIP/cBvD4MZk8vj/VcJv7mrehZSOKpBfS7QEhuw3YYVViNS38i/04C
DVPqctHnPXLoRjKNp89nvEjS1OdVIKJJbdSuJ5Mu/f8w/I0q6rXr3xaQxYbQtzxOFLxM97Rr6CWO
c1anIEXy85A37YFVaeDbWgKx8JBLa7YaJd8j32u/a6KbNSJXKcxsZLaVB/fW9De0mD8LKJ1/RbE0
uYaOrt98V2DKegIFDxsUqgTKRYi6z7XhdCn0sP1/CTumhA1JRcvFwQqlYVzSsroZvn2fXd5kjELe
C8KfeZydZP8knHzrOcIBPRDWn/Rb83Qbx11EGFTRJrChOdKqO+MPAGVTwXgg+EOHmZ92LvUqS3ZT
kN2hT1NU0SLbz0gBt9k0BeBfuny1v+uzOxku60hf7DEmE8Bh6x52wmFQ6iUaK2Zbfeu97hlN3yXo
wzCmWZP1/rg9NBm6Y8k3cAz6Ea6pQZGcG9J0B2uVwgfHHMUvM0/n6JmvKDoBxAX91NpBel4+xXGS
9JBkGKeIPAlvPepN9dZjItEG2JE02O6n7kD8rPtdpJk72pyOYKmZkrHaFtriOv2WVPmtFe1LD3YU
vFUDquWTF9VzvYnnHPiFsqUBLA3VjjGColYGwIYduwDmlRUwdFlJNQMReuhinSr/mUaw6RaaigtG
QbuZvaMDj7ve5PEPyfYSdCAs8Z6izTpQry5bldQA3Bad0l+ceEfKpU564O07piJ6C8hF4kW8jZhV
zMC34+04/6eTe7dfvDYKKk52GX6Sx02Wr80MwDYtCmFFGciGW33Ta6ncqv76JwfgejKDnOKKOb64
tEfhb5aMdow97bFby1oDJE4wTGRV/V3L1oDbwokdUJe2BGrVRfjbCMcU2xe0eV/meJnF4TCqBrrU
auZVeqi0eBJbvIpo/qfsZCacUsQJzVmsbTFDtkW1s+ajnnmdpwrSYg4X+cCN3hIoHQwskYa3Oq/C
RkqVdqgYtAkWwuTVklupGwcEZIyHRoYOmcjzI9Ts2P5WtWsCLLhGfZ3gRCAISPr7hohVw6c+xW4m
OvLkr6DSKKcyg+XscqbRu4MydrwqM9dQUHqfvY80odjqs8R+8hMbUEOnTNOqV/IoR/mMwe8xen8w
4p4ZByCg0FLZ4bNVybNkeTEquPLzbAqQ4TKQr79yjH00QB4Vx261k/ZCPgKMz4A4UA2Xhggfku0z
gD1aK5ifKjvQRs4LChxuw3kiEeV07W5o/9ayWetmTs5iTxro5wVLZGoRNQBRxdXh4PQHbOINDNut
vH3ZnrPoXWa/FXdz9W9rGaQB8hBgW+nAkQgGolOAb4r186yxfqxl+8tTDaQj9ksZzlLStDF9k0Qa
fJpEOhrde4NQfk5DDRKEgoB6sw/C2F5711CPWPt6iPHRKbzKekfi6DBrRc34X7xKnJC7n/DmKU4P
1MvX5TvUD+OZ9HTMOHt14A+/8NJwnpcNaEOK6tj0EqeNUUnFGzLh/yLRti2/BaPQh8iNt1KdJ6WF
Zb+VK4elt8wKj0jNI/LNZkUys33uNliLCQrdAJ3WsknvKa6HxLhhNwh7Wqq7AWibF3gpFIX/CYzt
xUSN/Kk1LIWAHVRgepawJybn2n938nZirh0uS7YqK3h+WtZpI71E8QsXsKmhIoOGN0R5ZEpgbhpg
OcD7ClPwZz8bY1YNDIU1NkEe5eK8llfq8hqAyMbqI4IZ0y0/JvWYS3xJ9SGCfmf/TkLiDV3FFas0
BoXdb6E5wd2ZOH5KjWREVYjSacwtRCPEbjehzTzf/RpgRNLzD47hLsk/JpQ3nLqufRyfRcXn3shj
rza9JRBBoYRK7Qs31H55cQEbIQ+G+vqZDn/lXaj7ANLGjvvBGsyOQIg3tF2+zbOAMBknuz//uafi
afiTDfy6cMna7i4tyJLyrpmM9Ms12P6aYXiP3PCMsd4gh6IN+qzCqJCuFaFfpPuHuUCDxxLQzRO9
GJdNBE/SumtQjDy50bwGRr1uaRakw4kI6djouLLg8TFzlq7ajEACyoJqrHuBAv3POv6K7mUi+msa
1evhjAOlT2UdTDlsrc71bKmMEayP7fbwm349tq0GhYwhsvtK1D2VtConGxcjw6fGRRuRpaNHU2M3
inZeDN/zKCnofR74r3X713doelNxVokAUQE525sk2M/ft/2BHZSXgawx1wkbRsm0KIZ+86q5LFwH
sASGiTj+blGATa+uhnYvjlzZepWPF2IpBhvFnTlZgcFlPVzwY14AFyB++1XIrGH3DiilXwKZps2m
Gxr/pGC6cuzCjuNCIUFX4oWFKL5xPv1ZoobTYgwYyjGCkpgvI7w1PaAyLkgkpNH0L2JsQlZoWqZ4
0AfPrWyIyBMclIC5jb5XMir5K9gJhgUFeSLT4gM68XTXFIzkpTc0xFYTSX6mFzFYHxqcyzmHkH1k
o3sx1ohVYmy4+nxj9NOekPWIXNUXVGw/csUzbTWXRNV8Fy2ieSHLjOlamQI5evnkC86/tHxAvDbM
h3mfgLjfJFJkTrz6T48HzWQyH1fxFUKqrLp4htydxfpgk/Vjpe8jy71/irJ5vjanx311D4KtKDMh
LUOkRFchAYdZ4UGFUAfUkY0HnQNI2nT+Chn1lNpTi51qV17UwvaEhdSdQg76aYHcC4vUXt3G1mcV
wRM50McWT+G6OjI9CbziYduEWD0nWuFJZ1hR1C7uw47LO1Dgrlc4sGwS+bC02jOW43E1IP/AZpA+
IfyvmQnB3XfqxWLT/9hZ2beGGhMqrl7hKMonjGRqhoaC43iNPNe+fTTkS5xJXpOv7KOW0y5MLtOL
nK6GGhWCX7VFGB3Z3fJnWugQsHDkoWvqUL88+eTWKPq5fpZffsAKkrGFvxrkbneewCGcJO3DgHtw
2YSIN/5LJWusiJj4dt00pmgdfj5ObfGiaKgQB8jZk4TaObuFbJq89twy9yyLl5uPrcr/l/EbDh9v
ueXmvhXnUI9fr3ZlB9wbxGNXJyQlidb0V3kgA5mosDVwcueFi5f5FcUAlarG7GFICAVtouwNjlij
Ngra6eLcQpfLBybEZWhlb+66vPr6hp7qKMhASx2fhSbuZMSuYznaf+InOsvhQHCfjF6d4rJd8Qtd
8uP48N7mfZy+oQjBhb7B4u0L+dRWSfRgQis/Kb8r8egr0zhydxtKvjWasGKN4jvt3/0jzITpsRKm
3A4TmZ4THpJvmbh7ydc2vi9IEyOJP5QZvQkZndKPjjMj4kcx7ZB8jUfuk5y2gdE/DvgWK5s9rU3W
AaNU2HrpbVepnPcP8/fD9yzWFQCtam4O0ojBWM9hJ6ezH1ndd06YEC5SGjc+IS1otzxNJq3RGgn9
r9EocD8yHt8owZfwz4ulUvkuEcFlbY0dLiQar295TFKHfRaSkd6KF8c9vM233uYqgnMsxmzRySCi
hXAGCTTlGYe3O+uyV3EuptC2Pk2MKlKnZj0cGJ2jCRl/bHxs058WL2F7zIX5WqDNRQMzCfkqcgY+
f8wczlFewaNLfsUtCJzwmSrRcMX1FD3OrZnze9E22zobmbfogtVAdEP0zteknEF5JNpPAPzTS0nx
Vx9LAN8wYhgzvd4LNYdd/xJF64ibgTwuhNbOpBuYBNDCWMCRfr5bpZFe3nETX92YKVnZ8RQeIbJ7
PhwBQj/R8UHJIRd/F7ziBjtqf8aap6URz25ZbLUXTS0068CucCLFXLMTA9VjtiLF1IOaEjYotrv0
5XR/0oiE1+/gznmiNMN2AVMeZp7NF0eHRy4iJKtTkYKwAyd9+zX2dQQBP+XLiUlJW/zWO/hN5pmV
FQThZFqpSpa4p3Hm5ezXRDziJNWX/tXRlcXiWas+zbGPPXo4XIN84zwHsjvfoJzapr+ojgA6SzB4
n/Ynm9nRV+dJB54kKjMa4ktEcfZOd1S8hurVUebHmlfgxGBZfszjrikl5RZbBX0s5jOwO3DMikWg
6RCq9/l2uVrvQaGfuX91XI/NIvWD26xz+G9IE3Yv/1DdZfIl4qtZJ/vksWDn33Vu+JjFP+rdhEYv
XZk1ebNqCBmEXARMZY9X5EBep1zRXHKSlsyPnqw7rOuEO6fch0RhiEL3GwOHZz4A4A5ATmagS6C8
Q57k4KQIMPTuHTt4jFgemCzkpMu9OwMbCTdlSdaxGaq7BUCyCJF8DOZGj2Lk/Xh6fF0srw08pIUy
MA5yCGCQEv3qf24+rvJiJlPT9uHjflaevfkMk/COKuAsbRooHJV4KnPCLYC8ZxBuVEJiNSG1+ruT
1kTQIFAQi23xZAo8pyDjINjWOg1YgEDSOVS0wRIiLss9KRpEwTlrqVBJDy1dCNc4J5QlqoYIwQFf
MfKPwgd8LrkWCwxpHu+829frAa8BzIVbNCuUptNfTQTDjKgqTIn/amxNGwEqo008nKsXrkCZYa2u
6tDg8ghFilfmYsU+pINhfe0UXY6HVJpVbbYPkW8VyKH1Ka+j3y/ZEHhe5Y8pKftOPsS4KbjA+qQv
XssBiBzg9q0CfiuO3b6EivEO3VCjYVlY0mYndwOtZu9ydaxj7JRfRg/hs6nW9cEj/1hchyaUzz66
Tee7JtBgbeZLnrWS1hOqQKqP18C9PrRExhPTbj7wja6cGQshswQIy8O+btfkzZwN+LTuDNUtaK/I
Os9NTxjcYEVi3tRb5dF7+yWHVHYchbbxPdCwNgiF0gC/t3lwzY6oGVvMb5oFf44rBeGJ7fxEES0Y
xLjM4n5fQhQun8xZs0ZsYW2tkKu/ZIDWw/rMvZ+b47XjRoBqWQq5eIAOG3MykA4MYVPx+pLkoSxP
jUAK6wjbir6qoBWI8eTO9QpvRz/1S7OchONHNnwOh3RfVwQvFgbKNmg4vmfqSP7UzzKbcz/UvbvX
+Rt4iBC2cRr8n95pCV8eXu6yhBtLP+VlPs3SzZa3pmwBZeN/jgpve6/9sR62gogBbzIO8Pq8tMts
Pu8EIF2ZXwquuSZomdA0KMhfX/DUV8iyS+GSCAAaJvGVRe6YW5/a2dGQamNtbxZF1XilvVl5cDAB
byIbkQG++dTmlEyTwNWSRmi+0EM7LBZ6ghqWzuCOaQGKyQB7AGzRhExKHwVDnXK1+a/yhX2wlO8N
F2InJm6ATFeyIO74tTUOXFc/ZvweKcyN0t2HOljnpxNxuwIgI3da1sEI7BIae9xUT5dce+8bVccC
kT433BJseGWnyH1YD43sB9zkEkwxCosFNZaTM8f6ep6ro2x7wod4C/0vQqcHndDbpIdF9DUbHgIZ
vaz/E7nwqH5vjgTJtPQOVaIHWPlhVd9UqY+SNixdwr4RW7nlZxfP2HJtXPn11kS45NUjF7bzVqCI
hqfJyE6Kc0nFtv0vzCLyDyh2i2IAsR1N+JmEkHy+HRMD8KMHStTujLFY4M/RBqo/yFJmUXIKcxNb
HVhYdEoW22PJ7YQemP0uLrbkjas513hHUFlkF8BtAB6OC1MQMUMcj3NSlnKfjC8dGQ1QdX4KyJk3
K0SsUUvkbM8nMhHArXPfDsXkj0DD+GsUYCLniq0giwu+N6fh7BLVA9xtTnryLaY2tjoRRG2R86UC
wORsMhxvaK5rzgYXpjyhyTW+mEtuOVQqyFLH5cWdpDBtnS8iztvHg8L+ffZ5KiiNFmb5DFFNygOd
ouLxiVM3rwRmO+kr9CFHZa2Ynbhf2gNwa09mbRbjfuzirqzDTZuirAIfsjCrmOjx9y3srwsguwja
As0csNmG7QZsDD8oqZoMC2ewWUffJ6g9oA5x73r0QkCWEXXth/+eLHXTt4J7BWjIFEc058b9uAcm
BlkDmNJN4tJ70A7UF/0ruQYfPsdzLavSCRuSpsQzzPpO0CD5XBvraKKNSqxmynpzWt1aAqqHPxCY
zvq16geEl4ez/cPICvhV+4+CSClN42sTzXGCRxm5T9RdrGQ05BFB5KNE5f02Tgv/vp14KUBaTxMu
8GDtgdUXsYYcFvyYBr6oi0SAojfjfd/mbTdeza9vxrv9QWHW2LCSW6EbXbxqgWJBhe1lTD6Ho3zs
RnRlmWJ2MhuC+bqWgUsADRCuvojjhFQp2GYZqrkI/lBvLwrXi35el1Sd0PVjAS9lHKdVbVV8HAzY
7p/3x1e6ga1Eh7jcwZ1bpb+aCWdlIsGrDNCKmp6Xeunv6n38nyKgDqtE4wC2sgB1tzRzXzSHUXR4
NSauVMNs1PoZRx+p7pBGm6/SEmrQYzWo3JrZM7EwmtqWxdPq4CEw/QGNN7se4e25CutMMOY1jukZ
rebvf3lzHAbq+TjZJckPip84BHGYjoPh3RBGrCX/m/z9zGQRc+AlsONicZsxbA92h1JbQ4KqYQI2
OKZpvvHI4TQW+51+gmyTt8Xy0k23Cso1yBF95Up1q+AQFD6F1KOJF1VyuHNL2xO65U4x2X4XHP8F
kcy6cW+5FpUuv6YUPDgEIBel4BP0JC0ze/c3grhVDzjmYK/8dwDaNdqa6kOJz30HzebjgU6e3WYN
y/HlqLskyBZDy4S5jA3o3tjzZBbYJkAQmE3kdlUFVJgQWmsL3WWQAId7aMSoCgqoVVLNTNvWQkGi
GuvCmgikudf6wADc7A7iublT4mJ8g498tILgY8D4RMQWVrXAtlmI0qvE3nGp5mFpajLA5cyVdycR
qpYr60yqdcGQ2VSa8cjdey6QPE6RfWTsh+ZDb0unjZglUD/eYQQPeJLmV1iYn9qnQ6yCFF9lmVvV
5cE9JJng0bB7n0o/0+JwoKj+MHAmxH7rPNtviynWQ7RfEUX9Fr4AM2p2K8ZMwuNi8vYmQrt4GsQ6
N4b9NQ27HkznVk0zzjJ0zIKuRVJWstSDWTNoCqpuns0QW/QQrjOm3B/EoYNCv2Dg32HcrBuuh+LM
7t7IL7Zsm4y+rAogElV3y0fQZ1fWkGP9iIrSLMmK/kEUbx2JnI8zxbxu4X8VZDbm0PUL/NsGO10H
TySiSLqUSz6Dc2UzgXFW3DgkGBBRGq2RubMP+E69XVBGQguSPk7wE38XR3JJ80DrZFobbV8oRVMa
LkVKLg8PQStKXPZ4d75CKNIypDL1qgURpgENx2XP0XP9UCO62vTUhZkAyQPvIyg0UxbwxQa2exfO
lCXsdyPZozAV9AB7ZQfYjmGXcYpMI1wuQwsfdvHNdFozia+w6G88JW07kSMv1CdKPRO4zoSPciRh
FycskfCLG5YPBcOlNgJ+ti3YrtkNlIMHeAlf+mKkp7nMDUWAEd+6+dRGS0VTKARrqB6PICO5W2kE
qf/m8qOYNgLEgtG2GSAKyKFxsY7M2AvfHPSK3ygvIPX4m7dFwwIomGl5dtUBejkn9Wf6S+LUUPx4
sfDEJ3niqIpXloG/2eZDFzziogNPUWQB9pMoXc1PlscGvV3x895DwS7MnR6yXmfQIivwwh9916EY
VImJ3BvBCwumt/6gBSdTzYBpboDIf1zR4B9sTn0pxKH87hsF/QP8p7WmS18TgDYRAcHLqPwqeGb0
aYQLw7LMrUlTia+EZdGx11X//W/K1OH6MOhV9bEQtdQVi1yMBCiiJWrsHDafTFXcBRhf6eUELc9R
l8CuH8X6NWuY6RCGxWYqT5VD3Qf7dcTy4Q+n80SFwiBE3e8mkNbZrQ5xLQ7/h6Ernqn/rZMmhOBB
DCda7LZABi5uWxTZ/qhDKbBN6ZFF+dDU9Gcs9Br2v0OPTwo0+SUAdB2BFt7cgDSufDSZmvgRnFAe
GOO0tK4oI9gMeDp4ic1Oylbdap/n/tpYcn1jNsS92Ziem1ndGiR/OdkrJgB9sCEQdSXJwTCfES95
abIDiqIVWjd6HZhIbPXgbPG4SY+ITyKSZh/xZNb5lF8qA3ivxUOzluygvc9qwT2A7E1TI+SgStLD
VR/w4YX/+TQ9GV/EQcVO6BiSVaiZbX+qzliaXyenSrS6dBzp47m+K3Yw0EmPXu5fHuFqhoqzMYVX
goDpECCM9blbHRkGfKbWym3bF9NDySeAGXNVErixshpk+BRnW4pZi9n1WmxdDTjaXlrpX6Z3TqwS
fPH4SeOASTXGC6oVnQTmm00Ehs/vOhwCAZqQCBKk9maE+3lquOLTtS6eQWihzF11lzi0COH9iE16
vy3AIPFZ1+marefXhMUyYM+p5NTGX+J3fhBrP7KuA/ilCYcZyxEUtdKZNgRT7XYPHnqr5hmZnZCv
DkkXQoG/vboKifAg6cOfVB7sOpZuEQnX1VUBKgKqXTTysJgkHRKGbbyPX/4quYJfSEP6H6sVFFyA
dGW3HrMhsYxMci4om1KTMp+jRJtxMhmOVIfHAN+RXTqP2uNd9Ql8u2yNYOMZqT8c/IWYFYDJYV4M
qobnQbD0JYvp2Np1XKTaxeUtrTjyWJ0HsIjowqdyRzgv0kRGv0I1QSgv4lMbythl01JmkkTBsacK
ptw1RE8tuW3/H6HP954PBpB7cw/gnLLAyIIn02u3kXYtF07lJBkYMCkOA0ZoVExb0n5WHAq5V7Ru
BS0LLAH9OhhdLbK4ErZQ/dZMpHn1ojUboHkuPva3pAXVwtc5zn2yjfZUUeYbYkrtYyefqnSZvUZf
3m51VTghjf86xBtnfLLGMCDeC36EiANT83vTAunkhUtHUM76997YTtYiyyjZyJGkWnZHut6P/eaB
67dw21t3PdUS4LAniduLX0Jm8c87RU3Ljn8yZlWKUV01TBwYtCCTAIoMyWrQgUv9oWZL7EPZv3X3
SxaDZ8Ot5YxCmBSoW0UCNC/beFPUCZdMehiAUTDHC+TRRUousr5IRBfBjpKG3sxd+MXmLjh0qQip
BHntardQQjFai2msWwcA20GAbHMjqWqeB+RHiPeoAK1cyUFSsSkTNXJfuyKlV7B6ytrxgirwQJkJ
pEOYTuysiXW1ypsFwKOrfAW1UgOoy+W+0w4WfQ0ENe3Gt+/QpdBnF8xwYAEyqrXHsuFsBaa6z5lb
00rZ/eIpafRdI6DGuuuhiT/pBo1Sgm3P74gJh3MpWf2Nv5B+tbF/SFTnpPj726fswFm/u3RUVt6I
tL2t2F5hvvK9Fozk/HsX/YWG83oL2cGeznENmStk3YGhZ5jMjkTfxsm/rd9QcZk45mB5yeSDiA9V
FwzEd4yyVML8gK3ryjKF65+PMh/Y7BYqy8rrGQ+HKMP3kWeL5TlMBK9dZ/p1HnvKdQrTEtHayTDz
HRxUxL4AP8TXcbSo4l1auNICKSzkDR8QShjelAyKYl+GOEJmmMG8wdK2safT3rdnyybJ8w8bK8di
YG2jol6DgHxoGB51uIifDgeZoX+daMVr/an7JGJJW6UPxbtJBIHjRzWTyQHfMT/+ktYXCzzfgPMp
2S8wxjz90LZBIQtKIm+fpuqYwO0UgprK4Y7lGTBuwwMHblDX3zj9lDGpwNlFpkQLuRh2wgbEThHJ
zCZtn7FnQ3pGlyDK1wL6jLIfwOuoDnu/wf7ZIrdWQ9h47F853rXjJ+mRX6HkzydwOThp56URS04Z
9QNcTXViYozmy8kpV2V41m9FnUD23vcY31kNLlgTIVzCNS0cO5+zE1FlrFgAD8TJO4Yu0zt6vLlT
jO++BphUa6FQcpkBWrw/97JldP2Apo3q0AkQW9syxKup/+gCxvaDPnMaELGE4ay6/EBdFFxDv2H9
q2rJIzRSi6JSr347micZpLd+qIIbDJD9PBmjMdhrWghH7PxIKy1ObD5yFYo39BTMtxVgE+fgcfQL
dd3WCnioKTTziGlMbjlwXgfp4uEb8tUSTZ8qAWBf7VLwvHJMRJd2C4hl7DvH7/w2ZejprT1AWVt5
qfJD/kw+RNQJtEuvNUGjiC4ioFfaYfDVXhVEBhr2EJPBmapdsHyHqGvbn0EiG30GMttyk39CsKPc
u0QWJbdp+VclOBjQ205E0tF6xxQ5IVm3NaeS75IPi7BEacY9F5ZZkdNBtuWHApz6RzdDPs///yrz
gyBPgX5IHMEKzhbJzzO9TrIMvenOp4q4nEsXfWeCAmmfgJw7DLwfnDPxRZOPB342A4FIrkV8K5Hv
6o+Lb6ktgdjaXSzmFnz4xkprWj9nlOFzKNYU0EhQz1Obtrs8Dhjjn3LRHBOXGvNEly3rD/J0EJov
D6MSJ58CMTVmhCEXHRbqVy+nt0TSRsS7UKrjj+TmwdIBrfC7rgZxaNYA1sy6Vk/AI3MnzZVd/7ag
hTFCl5LxcGBAlFsERiBqJAfpp3Me8LvqmIYxl4l13wWsFk3H3rZ5o1twA0+/R7eEhMRveGolp3yV
mpuA2BXW+7eZw8IOCIQDe4uSa0r7J/tsj7HSsvJVbwsCods6cqqhPCS2issmo24j5P1yiYWRDMht
bgCXp4kFkWVtAdm/UXFg/dfQJ5k2CCVrOnqAQhBLITom746QzwGjuQDm2wnu4urR4LYJIAC7P5Wc
AwWAioM6jn8bTbHZWeL4E0FHwXPR9xafInS7SZ097W7xVGjPNzhtBpSYjnYB+4sUfcdMRslQZ/E9
qwh+3q4mLyi/hJikuWTOI0LgqN2qPWNIBFJ70p0RVi8bqIjdlanqzsDR4UVIX6BRqdmaUd/0oNso
CD213NcFkj23+bRx0adbfwI6hn9nKiXQStl5ZImbaPlcQ/+dU+cXHjxFxlpDOu7XCjUiFs1Jfy3/
qusVZfIR+ze5urNRs8dxc/p5GYMSvEflLlcOQ2i6zbh7Ap6OVapqfalXJ4qitLUSQMJgxeIjcMYt
7Xb/Y+9TZ4kCmDVRZS0Bnmn3KPjO9DJb17cHOjxELSjsv3n0+R3RUrW4ijZPo/tFqzRlX+HcoPwt
PmvOIehIvwOLTq5YSZfL+phJbY/2UYsMU5yntuarKwazisGDTw5n1Ok0BoOedGaNc99Dl+5HBFlc
YYuiMJILsj8fVGKX/2suJGfbqqMN7okIe2WyhanfPxesoJq7Xmn023YzyPHNXFWTVcYve2IhiejV
AaBk43qrdS9FaJyGH/8rRVFwEg9WS8B//kjfIps+lAUwShVEkNsZTOnnaYybMo/YbVzyvOPqb1PT
74D/09mERHOyt7hOdleOkfQNJyMDkHVBk888DkLzSgynXXNwvZ010+Sp4xN0K+gEjwL+DIh1QQLJ
A8b9aK5nLFKP/e2ynZEovUwdMdLw4ZsGJ/K5CvZhW2ttme3DqklLQ76BS4mesDgcfbbpe2pEO41i
4fAWrwrAM1ORYm0EVnF24TobWtoRUOQINJxkNBnWDoKT5VyYNRQSUvMaqlaVPLEgL8d2RDm312m+
IN8BABYK0tqvFMlAHKNa0HutvarVTiH0YqPHiTG24wfqCwAyDA4QHZgIufMO/Lj9DG/M7mVPYheN
QSYCfWeKFPeU3wvRqpiUqurexpk/OSTaHkswudwvXhSfYMjG0O93LnB0lgVFAImQHBZoRqR+dFc2
eLaUFW0cqmP4+ZX/uG8KIOj0M14MFD//IviL/3pC41293UjNACj6KjVTYd5ZbTLNUmDz3p3oboW/
ADaBpHwnSdFHmMddDuLIbVh7IStm/RSDmauHgPmX3t2hGP9nDefd4U86VjTZom1hqxuyBrwXUTb9
PBnsmRf0fD6Zbbaz19rQYT9wJjySUcAFQGvBDCD4u5ioN1v0kecIcl4vof5Q76BtxlBdiySu1b8P
+vj/wDftQF+qrNGumH8KBgCpSwE/ClvE9L6UJFUhSp17RXNDBXpRBEA6yHx8GmGKxBsBovC+JOJp
mlk9A1ym2PaDg46b7cibzJ7Fl7CRBfblmDPEmx3TP0mS86xtARNSJ86xLI16xbsVI8ajP9FeDss5
HJPVFoP1BpFGI6ssutxqA6TTA3nqaT2IRwgNpRN6RS8/6Z7c/UwV0wc9QH9JDfWWbTp4jySr49TU
Hm+f+vJYIrsSaGXZw4IHO/n6DFYNL47oN/YCFKSxXHKgpYiHDyfWWI0aeICBVpRNGECW1pM9TYcv
Uf4dEllvBg/LxEgK6wxQOBlbFz3LCgHbfExe5KmkklsO5MI4qIjtfCzbLtmpNcEdEPclfd+JgiaU
nsUk70aDJZG5k/lHKsBfC7JgCyjr2ZkT9bBgUTJymM37CFmRBI5Bn5VL57juFcIu1lpyrWK2yTdT
+mO7iCqCQ/eaV42q8rP4DXszZTRfq9a1qYNmRFQh2zdmunjZ4BsjshFWBSH77d1x/p/9uMN5Yo6Q
ejLwQ6kIDIPCY8y+cR9+fl0Gus0iEf/zh35xhpW1zlapyR3xnhPZoiAxRI9ntA8+ULsk/x961OdH
S1VkM/W/JxuLfFWp3gsVj1tRiwiUU8vIVa6i5OAyU+pD3Dja+bpdXnZQ4Rm9KvC7er+uEBoSVpeC
/yoMqb3yznF9GpML7FBAOAziRA0zON3eoAxPucHoih3XGvkCHsttmnudz4xwgJieQA0hPHEq5Bgu
jHbSUcQE0B/htvYLwJYUPM1YsVeeQ9zGhqfyBK3rBKoTyS14q6BAjinma6yLf4Qpq2z6RFXj67hC
8Bel1KM5WRIc+djX5FKoSP0OpVQOS4wbJrTzgjAZJD10srLOTcSAnOPiKgQ8qyplMV/+MlUgaBO/
TFOo6EqhBnwjU4L2hrG/4BgsOCjLc23zGhS8zpNYLb+AGkTPNXGXNjppQo2IRP1nXxG0fT7Nt3jG
TptS5J+LRlSRgZN7iZTCWFQm0olIFE+bMQ4++B6SKRHqKdMJb8p3SbvE47S47BVvX+q0s6h98Fv8
DxSb7+DBjj36NshtyyRDEnofYnm48kDEirWHN/0TMMn57i7/mKAPF1V6VPvbxso4tQdYwQNpcl+F
XhGtwKu7KnmJTGH5m/GCkWtC9Q5vomJ+a04pwVFqN39BpE9Ee01MZX4Ljw20+AxDVdz2qzXEGgNN
9p86N6s0l/k4vOPpFuWoMyju1YSA4Ad6YHLXpgHYsfWAM14mE9O1uT4PxLVHuLYUtvzV32gTMDG7
ksjKaQOaPcvc/BvjKbV7VmDLexqlFCnpU7YgpF/XKb0yV5L3VYMppDg/nxs9tX+r0p4GEW5+riea
5cbbFUyvL4+fGGGA6NX/kbzeTLJJ21Xj6gymlOsXH2wOUuejuIifwfAC4Yc6zM1xnY2apgtnZtKc
PkU7liJpeiYX47ddHnK6YwK4boii+5fJDv/jEzJXPsdiX9ixlWyWGt8jSDSlUOmYkcUww+sW9wJj
XnIafg7ci9DNdzOU4PrNr1aZSQ2XD6lr6uATluD+9qckc+hZobx/5B4HagZm81KdrNUKcakP2K9s
z1c2ZCY9SVjB1QQkOUX6OKzNTc4QlUjCJh5Pk1h4KGTqzCMUoJDmGSt1bWWCOEsJ64mkqisBFWNW
7mFNTkByjddkI9Fj+5oa/G/Hk+qCOVX75HisnvA9UJOP+fRAfDEx4JONRToRqVk+RLRKQ7RcF1F/
rTLl+8w5LHv0q6dFxfolxXs7rgbiGowvFa62acXKqlV/J/LH0tQV8j5swSN1F/Cifrj/pDQEwKT6
7u7gkdbsx05xuituKJXuRw+b837mKemGi02bJO/QNsvwl0QPCeGDWFebg45hWQlUblhLEvdAO8QL
jTFmFaMmadjQrpB2pR4iEUiA8q5UzpURWCJDU/HuCdUhPAIKEjg2gtO6Xu4fj/rUipWzVEUHY6FT
B2Od/yatCBfx+ME1mBUR8HLeaGlECHudLuL4f1orc/5bTJ0dR1fkEAIud7GIy5ikHOExD6ohla/4
rewvIN2nSIL5C0chQobXKqVr49AhzUZa+nljoHtBPfS9X0RonVGU+yVQCEg9E3/fS6v6bijNnJ13
FHeZ8SYrduquAHXGJe9QWfb2xT3uy5IjZ9cTyBwijuz5+EDUFTQ2Li4+9vU6lB1VUwdSzRLc6sU8
nbzGOIw+iwABJLGPJU9RLkdQmu9/NfsjHweBje2LNvf5Age6Xuo5EypCbSWafJknB42II+KxI7HB
LiuUZa80SqVTDNyTG7etk573YYDzrLnd5Zx0UMtArA+sBVv/Fyj/TpY0hJMaaMM3k7qYJrHiskRz
r/ugpEn1EhSHpsf/FYAcYWV0ZbTvq9iCa0imiG0O3RBUp6jLxQA7kYoUjL8kF/ZxCr8LQXS1ZXcb
OCLe4Argxr87drMBYK84zP/PntW6d0xgcKngS7lbOskYSUw30Goin6PPMzgVnPS/AoDBMJeMnO7/
AhxizNbnx1t58li7BeOgO2Aox46W/WpzCa/Z0ySanAjfUGoAlhHpXE9TqPJSOPZwWr8Lrk5cH6LX
fySFCkSmeRVXvPVMITrhNRTHCxdwcCvOCpXzzZ5ndGeuy87KGjtsRT1hOxOAPDDS+gruudXPv2BK
FSAH2pKg+A+zanOwTXYwiEcMerRrnc8QCosmtZ3C6NEYReV8eEnJ1dMgpYH58y/YeiTnzhZYp9zQ
izGLvM3wjISYp4v6wAsFYyZNvp6Qb54LK1rUj0SzK3NFvUP7fTqEeSpM9lyP5wHCyZzCnujdjuBY
N265aA0+H+ygNvSPMjwQNRfvxsTsrVdmp0x7na6dHUWHg/1N+N/Y7IqjSQMSUGGbtPrnwWD4fuOW
H54PjM07Iw8PTXrCaBtVSz3krznONvbyw5UjLWQaX4Gok9jkfJmyia3HS2gXCFq1UvEv4aJX9TNO
YmLnW7z1UKyTEKiTj57uI4b7MNz6W8SEP2Wy9xiAwkl15xzne+6BIIpzSMR0jGz1cc+mrqltY0zj
c2qRifOnq/LXK0Qq9WvJ6bCq6J8c4kiDAh1w5UDHNqJqhRRxhZCRjutvB24BUblgfVwR0iobSFWD
E4UFeDjgbkwVm7LzVek+myDRyLcS4rKYdaJrrFAC2PTGWf4C+9LyLPtHerzwrGVFOlrZ4FqgxqgW
yhANTJaS22KWX0vysCKo+PE85eTS2W8v6/wecOiiuA2EjnZ8ZaU7US/0Kw7S/HNCSxbF5iBUjD0j
aBEM7a4QazQDMoiLNnbuEHaRVeTwLrTwLS1TloEZwhhlOZBo5wMJ1SgyxShISovAvhjAOdGPlnVS
9VCOKDUfJMpfnopsTg/KtjBcB4S60bxzUGnqrQiDeokhWqgzRCHayFDdH1a5hvjxpBI+w/+vBg78
KdAa+bf4LfWnxC5EsFDSoBRKFlzvZk7qljEWZFxAXR33PyI02RGRrlKiYtw1og7Sg8Z+zcgLB2sh
WNR06M2DPyX/fWzvFolHSKLFfHtgZYCtiasvY2wllOM2KQGVxm40dqFZFDAzWezNPuk7Xz39rqw8
HiukwJnmtoUchbGCdT38GFHq/SwXmUOiisCs8tA8jGLuapO/qRcdxOD58WepuduFpVD7SpU/Z9IB
rXBIM1EcbFYN6GxlzkfnpHy+M88Nh3eFTjPWn9zOO06TyGYnznsClRUrNv63y10j9Hhc+0k9a9nx
EU/aI/Et8IZaF1N6M+MDL89tSeU24DEcgNcoKUilgUKr4uFBwVCrdaHKpTTOPsPHowhpisBo2ImV
kwhhDL6+mPbbUeEjnhR//OvHn450zxtNsHu5OqHTTzq7CVV4PnE6lzWuwPaBAKX2l7FEU2sfukBg
VX4tk/Dje9hH0mR8+4cOEI9g9J3S3B+LshthHNYu2gblj8Bc1hmNZRjPPMDifXOffng4+AOZXuas
r8w6CGCDtGyc4en8NrlyPUylu3vRejuMqyueYAhpe4F0FMY5FnDrOt/ImMstmhGJK3Mtcn99AWvp
+jKmBouhxiZ4pD8B8Up0WMtGVgL/eUxah7vVt0TxbIbGRG3wmatPfYxbRYZZNW1hvYiiV3qofWS4
qzBg8cxvJYD/F+BHV+t232QVuI3eaV6IUAAy/Zb6O5sPFSdM86oHc2vLaX8chTtKVyDI3wbah6Dw
2cITWjq95SiHhn2WdttOtTMdmvsvm46lXraW1SVN4xdD2jI6mG9inrsEy8Ql8cPAQbi4VG8TTNoj
EydQbC6ODmiCOD7LlCKfiI0DIt4Q9vJvRrWVhbNc2oRuZCu3cBnEdIj79TLQQrilAj32/btqcbdW
hNOToXIcPMJoPBr1SMHhS5/8Ky0qSSNAU8t8fQswSo0oVGPe3UwpalbkPLNwCs7uKo5TIGdX213u
jBlTmrpDfp56x1vQu04R4hXWapi25O1MakSjyZoOtK9UW4pLjYfo5XZWFQ3LYYwTqWZpYrKIR6OP
uCcfjbx2AfExp3W4mvNDWLtkOCEyPYbvt5UrRkziLeXgUvrWWb7RYNB6f4UIXsPShplJrfwGC4gz
h1lKT+Y+EW9e+itHXSCfcGztPkHC0Xjq4HFFXwSaqpFj3fkgRf6oUc7PIaP6IXIFP5l5zD4mjI3X
i6OYoCukK1gaTzi08eVtRRNmAJohQ3p5sZf4+dwRwhGrxns1lz9QE98b5GZpUGAokIBcEEvra+EL
n5YN+2zc9TX7d/f+x5WUMvegMxKkuYcWyaHxyVixBLcrWSQXm2qpUSX2diJx9AYNeqGfKLDntjuF
W2G3N5HNmYc0J3/qB2FwvFwOthjw90ooMM93fZaFRBJ0zQdvLOZcXaYZAje6tCmtGcGZfol3pjG6
Iu90Qoj532CTqSt8RjR6WAPWQ+zUOV3UNcWagUGIze141VYcLbtIIEhtHvUxChvdHZicswxDFUsk
+uY7I0SL2F+WhyowNcWqKmQodD6mG0JlnoQQxZUodjJDqF90ja0nWL4rBNmJOdMig736+3yDzDkO
BadQPKj8fUaR1+3GW76kn1AF/Cq4xYGN2bKcZ/bYfm7ClU4YPgIIV/8q19bjr/0vzlXy3o3+yTVS
dl1CCFL1d5ElQdd/XB/gjjBVEEpqxIGPxbLwGmC6gZfeyAof5/+6KCTXdPGtF8qcBH4n/dRwC72C
axGlW5P0Izl8S8OxOsgJ4h/iG7qNM+T70P+fEAhk7439Cn9kSH/5YE9YVRhv/Il/qNw0r/YvOvEF
4XQMyuX7gRR+5wZuTxR+9PYDkr23Pn3BgWdTiA64Xi6IrB4g39gT7dHoxdKkjHWzgSj0bjTsagZx
ld7u6ZWKgK3b/7EynwP/NhoARXJ2hzGCgJYG7gWOTphQ4M4E4amZjYlB0PZdikjEhZaf+tLNZLnB
NkMkjmnm+BnIB7lOe3tG1GghZBi2BRQV4iw/PdaHX1LN1zdYKfVGwXfG/bn9q+8DaqHGkbpdXq9o
4nzYL6V2thwWcLBgklETFwJwc1+cu5pDYZY0U0yJY8TnIHSrZZQOF2ii/S5p8zNxdn2iNoIp/QPf
HRQfSiEP04Otv64ulTBRtdzI6HyHYGWJ+mVEV3nNW9eqYVmK+86qD6LtM2bkI+XYianyElSVJMNl
oOssVgOdE2cR1yXQrXE1uv+ENIjCcHoa/+W7fLH3kB+B8BDJIwxTiaoxsyOrXelv9WGEx1xD/192
jyVNI2K01aMn6irB7ZDhhwmTR0FRriyFV7mjy+5uCKYN6yEZJCw2xa/8kPBkHnLH8uRGw59vqcuV
GEOzY7+k6OMWhVW0r1ngKP29fe2BI8mHxr9EVNmLqzxsFPTTuJp/knjlv8US43Td3KAz2Y4HnQi6
MkLaPTC/wjd/SPrK+9n7YBm1A7Hj78Lc4A8n2Xs1x6fSum1grkAVtYTJnXe16mmnLDLE41hIPNBY
HPaSHHxTXNwHu3UHn/7E3eR15EFz+agszXrRG41EunN4g7mnai39vzFCQrVoX8P6DtylYWMudjI5
VxwVArRPbEZtu14hyEKzSGiv9fK09ZLPkJon+LE4+WgsKBF1+e7yXmNEMTdGbzR5pnV7TQ6a6oNe
KKoQNfrE+IWcbCzPiN1G6FSkDF8wK51BpupKFw473FdL7jIS3OKEMqmL1ogvYOCQb1ZTsNoVQSHU
68BYM+k5rZ9ZhNvi3/vX28QuwWuvzExrTGU/YVXXI5YSgQH5l4XBbUfvBEKfkrnjNU00s6oBsr0m
I6573xVadZNqIaHxuYCIV9l6mkgr5S6bsZpr/e6H3lnNTT2ObAsg/J90N2pucJb/TpwprOSWau9C
N4BuRXL+3p3pcu7cE1bhDm6Cm0ZfgLMNRXVbcBkTmlqt9y0c7eD4vYEXxspEcsiYw5cPGLFqNswh
SlNgTDn0Vh5sU+mfl9CTJFGWyeBgCTemFszMEsTPvITcFZgfMkIJsFEOlM61WOXweE/pHpJwGy/I
yVRtnK7EopgKoNGGwFYmjba6XQyog6DQN9+PjKeF0iibHwhIm4xHum4jzuVGNc13UYGIx+ldvadP
8zBzsW/jCJGo4+7Zsf+/A1VYwi7tn7EOr51Z5/N7L7Vsv5S5RFQT6RA319wYh2OVxYiUuo/n6CYM
H0WBKtWaLjlDuhtGwyn4rPPz2VindHGMb2VyGAmHEJBVhltw2DCbRjLn7GH629m66pLGBiuQUkmT
2wUQhDJaQQM2UyH/m3EljLjH1Iu/Q/JiYgn54YbAW1pirzgW1nnGVbQmtYcaMcVHe3iFTmGs0tfH
CRhB47EY8nm+idaqBnVtl7Sdmz+3SAPhq9OeaxKeFdbHhYNrtcWKqcAbQCL7BZlBgN1JsBQ3gBbo
sH8z35nDAgZTAh5qudPdfpluwczEb5dyL5663azfIkIhuw7TfPxetyMxvGO2J43WajmMT0dozv8e
PVOyUuPbkHzmAaiT1psTRa0vBDVCydb2xNNZQMTYu4Q5+8C2QQSZo53RXHs7rJBq54tE/9CaJnUc
fkQNgEnMteG6Dng1Q/n9FkpB8jruykBivVdnsuIAoGA279s6tkvd/W695TCbkoTiJhN5nNpxA8Iu
3oo1ziRprpLI/c35Im/mnvsonZB9qvAlgFKdITLoGG3PwXWmLN7yL28rr7g8PmVU5GywU4vGjrSS
Y8r9HmrJhjNSn43hxXvViCaQWhGXjIRG1iHkIrQt8U6q4KpIpHDgFdRQQ3/jVyQAgaLEMGf0MG90
rPByn7VwTUx2bp4d2Uwiq3qMgN3hnbgJdBDF839/W0enbulU8+l2r9NrTL7kkCFm7YPZSyELYmoq
N/p4bDul3/1FD2NVkSUs19GMjLHIrQaio2+GifMtHP0NTeQrw0yLSecX+LZZLmNbzmfWTwLQTSR8
RkJEhzQ+NOnslaJozrakpLoy3eWt0+0LPffMkUsR/iggRAQPexU8prf03CB8oebsKMt5v7U/0sPw
dUmCeX+Irh26UR+CJuAfFtwOVfzIyADUfTXHwijCS11SGSMMnlnz66hMXOrm187kwl140UboeAjd
fpaTFG5xsPJEUV2KApEWB3yMa8sMj0N0fQ4zgYzdxTHqTNqEWlGFy89GMsRXaQGkJ5t0ow9ZAYFF
UhC8TQLQ8ZNYBmjFldeWWjqdz6HDku1YFwv0aGl+FXHQPunj7C5PdnJRS31FNaNSkFmFcUF3jGJa
0aMh8wAylfambHC1SZZaAQeNPbJCAawy4IGLRcCOI2pZ/z4FUBFMwLajD2VljJJaDHnWuqze6qLe
o18SB6CpCkf3FMMNFu4i0kRnfb3wgQt2h68HckeChX9+qD5CHmQNFkZenokrvaWWrAht/yt+Pyb0
obSAYuD48DtFpmeZP1hH9QKiK33f1DDvJBYboyZ+PcSofLGP0LtXktazemCekiNjwVvwBaT5e7VB
Zc7FnqFczuHPCY716ehvfjGT+gymjWPRaBmMTFWWp8TwVLZp2oKiO/lcTg1yLhonujv2BIbaBxbC
7eqMbUXZww818Z6PGsN4a/msujVRaMX9PiJRNxWH2HM1yR0tK9q/eqGo2yfdAbTCcIGc2FSDxZ4X
bOFd2GY86bhuhxHZW4BTAKVFYEHhNOqfjct6wQxcMU/6KF8p2cNiGl4fulU6viHZ5TgodUlLic1Y
kbW5/U50JF0zXho0ASmG6jRbfmQ06y5t6g+5T6B5rpMxcytdeRWE6Y+Ei+T4YE34ia6p89e/zSTH
RRms+4xXgepNX6KaCTZK4t1sqcqgvJpO3lG2vH/4ohLHcCgPuG2fFl8HT6RdhUhZv0vDZHui3UIM
6f+3kfTdV1RXYc0rzd6plBTWpFDtL6JOImRobY3g16G5wM34u+n5GVWRfqEne/R/deFTiEy9o4MP
FRtSx8Hvc2MRxSqOIuZaatW2TWmobqeh+wU1MR6x3/rvoRGphwdKJECzQT9GsF7V74jRDuOVZCrL
dEsGDOXwaJVJy5r0MDtZUntzcgH/KgfI3CfNQFJkzlCOnLvFla7gSTORKM5euj3Qly06FoNk4a7a
eTqGFratqpK3r3kghMXI2BvWrCd1E0VcJ6GxnXTeAwoRzC9v3/+dkKkVPdF7+doHMxYXQfWMaSdF
zn4zY1ELCA7wYupaARG9R+ra7Hcgahl1RdJusbMN3vnJQ437Db80XtUQpFMHl/oeO0QVohcUWDcR
htiNQqGEN0pagXriE+t2px0TyMFSF95ZXm+QhZiWXOyOffM4fZv8ZW9SWp7V1joXDfGqh/mOUGti
t9n5/LuvnPchHog6dBZFXUrmtJjYKU+dqIl/YgIfzDb5jq71Nv/oy2i0Rs6VCK5TCOhzOReJznku
oSmkZWF7hNLS9Ck77hNZ31zmlCN0WDb0b1MMieSvdRWDzkALDEIKjGinh/f9PMqJriUQrkpTXt1V
o4oZJB57EYHFgESNGaWZdwksrdtEMvmG3l+4GkJ0TYgLf7Tp08B11802egYA7SiFy41QcHasTeF5
PzWWGwhY3EKL6qcADuzNSFjVwAmbVEPeHu7vRSH9r44FNRKYo2QB3cvLdSi280M0mdmVzInlzpgR
uNjQ4D6+lw+WuMRer7YpW4rPHj+gWNXIPz92fRfZh5ItEuUNHecndm7Gqu2gaXsdjWQfYWOf9TwX
zxaRWxVkRyJ/qQxDRE92ohLJ83+ODbCsU+5XkBTIgrUnpI+nSzN6/u/3kF+V90xWVEuCi4aiCsmk
hoPuN8vKtETda0tS9M0Qc7Iz/+4+xbXHyzCYsrBDUJjQKRH9mfFNQr1O/xWzzhi0Fiu4u/buLcsY
JqnW2E9C/HW0JvXzJJVuKXbJwZpVFGvBSRbptZapuOnOVZwj5AcFSQDwaziZ/hD5zB3dVTjDaaLn
L7NtCZ2zsqE29vzEgeSX//VnYE+Red501n+HBJSTSo69nPT1YdK/KJucm9FqYyZGxMryDTT6Clzs
TjtV6EQopUp5Z0lfD4zfWIcD5LyUUPh/cijQK9r8idqUE8dGp9vdoU61uqI/VupSatACiByU76kQ
Mdf5bzyo3Hf6XUbHfwdILHIxDzUkvBwdNUUDgkFoIrPjZO2o+JUqxjEZQF+4zctEB4uvek1ivT8m
6AKT1Ro493Uew1dhZc71wmjWk1GxkG16/ytJjDZ2p6bCoNyLsxeLuMFVfuQGCiOLcW4c05sYGKiR
0gGaMf9/hnB9RjHXzvzNtUoh6x7ZqbuEskB7ZtUKDkWi2iRwAahwhcEoc+toeIEW8NXzW76fPtqy
4F1F7VuFLRaT5stsMWTsbV8LX8wKlJYBleCdzIal6hRkWLea5Zh6Sv9VNshzFk+gtVbxq0LnKfCr
aiDbFgpVLg+OmZiz3H77Gde9QCNtLtqlO0Ef3RcPOJDuCmq9+JhLwupQPhT8bHyYostwoMjM/ZMg
ENccOdcmPIIV5ZOUAkp1KjVxd+8cTPy4oZX49XR4p0Ue37ui21Gfy9g7lsSmOzBiJDdKTi9R+Dfe
qMvyjDO/t2PJ+TwqvMmr20dDTjOR8jv9k5YjH5+qzdz3zb2SDpNe+YkAaNyziDJEhgnzbtqFtKCD
pKINDUQ4oLVsxDtYfYq6VFofFZEzONd9mypcIUmoye85IoOjdZ9hkGMie+BkN3YLvTpbnztu2eFp
UGXRJAyrCeVZngiLB1KIzgF9Tv59dW7bsCoyV80lOC0zASr0EuiaYOlTzEhpIL6CVlBSNDjG6H3d
d6ekx3htyA7KWuY14VIYDk6V9z510q7UvTcPPEMIfwNUPXNvXbVaRP65dEAhm9C9UaR67eOUgAZD
Ja28eXKi0pjvf6Mhr+CzIAUGPN15gj3SpEHIjcqL0OILCudowFxz/u2UnWNcAlYckNsSUoTrzX4D
alWU6DiaRKM3Z43hcvrxOoQsbg116tzowCzgCyVh6WKtcLjhCxSDwY2Mq6ioh2EhuUHufv6OjSHV
YpoVILB6ZQ6q7dvgl4Xt7wz1zev4t4drL9SnZ+ZncEkXeXfBDKPg9jIuiANDtTdBelk4PmwPZk/P
2Qs8gDBklTORt/clhayZ8+8mhnYitm9XdQJoCX0HwoQynpB8ydafk1DmfWYaetoCxo9d/8YTM02V
CP6PkRuq69USuBnBSykRc8flSY3a07IvcCPZlfeYiX+jq7w3toBVPxFqVULCVtSaadJMxT14M5Wy
FpJ2QaZ33L+SUntQLFHonogxfptX4XDpUJkdSfEABAA210kwKpUPCDPGi0I+v8CwryMR+Lzx4tfC
1SaDtVLpt58wPWKo9DNtJcaRvRQm4YzPhuxvnvjBLSDixK6P+aURapQ8KvyNl6wY6wy2bpKFbPn4
iY4j2R9jcSvABvv5/QV491tkwER/aGIcP84egVtQb0Mo6vDTyAFL+J/+6QwfmvAez7mONPjrjpW0
E+pkOMm7gt+JeG5BxdXoIBidIVcFJ6Q3ktKccCR/A5CTFtbqU/xpnXKLsKXLdNsi8KgJTKdAex6+
pJK6IKMsuaxlPrB1eNYVzitPUv95cEp3SHesCzoXC6YQJNogHdFDwSg9lDjHoeK1mWwdNdx76by/
v8AviiadV4GAe71jmYIxIY3aGnOqpwJfyKymh9AESTTLiUHPrP2BtXrbakOIb1z/ATRt2Bx3m2uO
E4+OGS0BBFTubeTcIPptfPBDaUFsUB12CFPkfcY+HFB3NqxqCRUWXV9mRixCaLIoneuupXgs5SVF
YOvojy0qCR1kkXzrm35Itc07lkv6zbKcdHNJl0x3HH3LQMWTWoQO5RPDXSTvgwbKo5j4GFkEgbUf
zBmtL8m00H/ufAjSkea/tBg7j+0BYhwVyGHm2X+SfEc1RmbyzmEJoN4QORZyyRlRjPwpU1z2HyGU
2G7thGgDAdnGBnjhg/vWaT/0swXfiWkpHzHbABrBV+dmNUcI4KN+RlA6xIGNaBbkPsO1l4b4oniX
d7zGgJWEfps0IJ6tfvxVfVcpFCXjB16tL31JU9wGF0p165xABBdO7zEmD7m7rrJ940b7rH1p7uG8
VatyavND54ios5+F7nyZBjquxCRMeQXHRGCJbI8Q2eIrnUfa5zorL0KMr6V3SIP9ketqokmGyqIB
31/B98Tvp6BGwXt61BZarp7CtzjegcwS/bDmCP0e4dJteTDBxNUf5uHxSBxZzQGh4tcsgabNVtw9
Q9CtK2xGi+wJE0AnEwxLx7m8YlNpEN+viJq4UeNFMbRsEJ54qNK/WsfZgt6n81PE+2nyENUp9I0A
RMNYNNINc011VIEUApQNdlCQUnSXcJsxDihdaRK2WshfFaqYlwN6H+jmNLxWTduVjI85X8Gnw2z7
g4WkL3TDL9rS50p5Y29qd8LFItswxdBgRmy8U+xC8QM393VncGdywcJdEaGcKN01Y55xj6MJFwKq
kb75TFaaij/wmFxhcTXNWADSBfptZo3TgCl/RsjDnuPAAkSsw6QhMfm7nPf6yNr/XFqj0c1jjB/N
s/1zqMsmQmyoTu0NCKjIQfae525iYijUgJpHtFkitKjwzfjR7jbz698uA0UL7YwTTia1w0mxNYiN
PeVBbgzAZwi58FfpjAGhtELP4kn2qVo0eGcQKdoqlZREGbhBQLfJr9cZowcvlhDytdgOytLUXNZG
uGW8nppwHNVcX+mz2oNZDga3KWztM+561hYqzcbm6RJxIafvbfsv0MHghqMqhn4CzLq2P1LMhm/O
QqcP5G0we0qHaNV20X2/u7JvfqzCPbEGR0gV3xkr0efzPgY7u9t+pjvKoG4Z1w4k17mnpfPz1728
JvQ/bIMU0FG8GC6lCBs1tTNb87X3aJA9z2GLvYKe29K2PLYizcTX490a+dpF7RapIMmN5M5GDr8v
rEZlN5iEOudywQ1J1kA80qBragEshzCcMGpKTg+FHLW9u8ZFM4ILO6LKw+6xS+SA1z9wENQgDDWI
iuJpDrw7T7C2E8FN6MKDGbG1fKSjpjxzXUwxobyoy3fAI47gNCgsJOeF1fw9fY7gTJjZoJPaZE6g
kKFPh/J6Kkmf4FIPNue3fMOdZeLOgqCRKg/LKYTVQt0gquejyD2ukDDDbUDjNLwmXoFhI4KGV5XS
lxSutvRt5XhPWapyKkTeegT5GKZo7SAOl8Kdw56fQHsf9cRI7NjXF+9/jK0ujmzuB2r3I3H6TZTJ
w6s4w/U8NPyPUYuuFVLBUI2hc+3/AaLFuyKmAlMhfIrKGVRz0rxjy+bEhFLOg3LF7/LWJZJZg+0v
bi9DkMMkXZ64rT3/eGDlIsgci6qr2i84sbfnJqy5vIQ2r2IcUZM4YMy5YfkWpoLvRHEizhbnXg54
H/FoEMWuLfTjPeGmGpPLHuW/14+XzWDiaGoL0SYs9gNJ7KUHZc8JaH9ykn6SJ+Hif9jhauxp88lx
Dz3IQjwWFENGw4jf1jeWGy/iwrSAVBSV7CrG651EsLpmxqDG+WtZV8ZNGUx8OjoAx6rm/68sRar1
azvRgwt0DwlS3M+tmbAsfeoxNhF8e8vzafseNpPqnaJFcnYb02exQ3ez63wkxetCh7gT7144OmUv
oJNO8hdAFnmHIBRG6VqE2xeKYvFS54EOaEN+H2L6I/JYMEn5bATUIf+WFVtw4P8F++ojZli9JFxz
ZdealDbhQp/3c8ax4nzFcHLgoNdjVN2ED0PhD4cxUFxeorxCX5vFEEUJP7jJo63qlfpNwMqM1R1X
l7jgYv/TMP2QFbk3GvnGeaXCk8ktG5VlpCSQUHk1xL+b7NwdLT2xVRfNEOVn2ISf/nlUk5rDBZy/
o3TNSkirLcpPHSC54Y8pp94VHe111vYhgbgxmTVNgqoSyTfNSSYUh859PRqvIjxtrUH19pdm7ljQ
pYbAdlhMT8XB+rZ7cLt1/x3Q700iJ9PZldPK/NRQLke9Puzwhv0kNC1Z58K7ymoo2Hkkd+vpj8Yj
pQt0W3ue3qBzoACI/FyXTtQAjBetEPQATc/R2au/LkdkVu+40j1ysqIO/lYkzzAmzdRbAWavEg7g
ySZNWIuQGDAwvBYY8oQu2ZZ2tufmd9iTWJN7om7ElwW4c3+p6FlyELA9kiWiiDYU2u9iEEmMzeVY
t4qs4UeurgLSkvvY27wSU1g3HRUK3qY5Q8C5CuVXjwqPUvst5ZPVab6Jre57Oh7VOB9fIh5YpXth
MqgBSWmIdsJS2THKTrhbklvWrfYNRGrKszYpbzm/Plu9e4JPDrQdbxoQLriQnPXXq2XXH4VZW5HM
FBW1C8ppW59YIs43lYCB3HEe2JbCUpdTn9F5hm19fjlDpg2gi3hObd4z/QpGECjdRDR9IuSBcO5M
wNTnkU8jqrJjqlLRtqpq6sjwrC1aIhbVaTFPbqWtWC/sDs5C8XLvQgK97TDa0mKKc1gWIUof8wX3
YPnjXQ2DQgbn8MAFrmaYP+ihuQsOyIb/i+SzkyCQK7g9oNiGxz//nUmmN7VG52ef2U1O6H7kKfyQ
G8CenpWqUI+TwC6VUHUJMeCgGvAglkCcNMs2ZKb04bUTjUnEfpv5hr+t1N1ETn6ZOejBKqtUIZEC
n3prSu/jO6xU5Ol0iw7Sn3ERzPvCKTidUVZ/kNGiNeSZZGwDuAkHdaq4Onxd2V4P9Mc//NOQcbEJ
QoqgaJiUcCjrLroLf6a5geAI+D9/sEMqwhmv+91b4kW5LXzX4cKssn1j9yFPDCB572kPW98gyF37
C0KKLJhRJJPMjOzFMoSp1oDvVNZs1COwfiZuZB8ndgHgumkDXBq4OJDj6IJhDAIQUvcCZeZjn47X
okx0pErvPly+vy210/39o5pQFQYnVIy03SVGfCfi1aqt1IefGa5vqOHJjI8N5w/HdoIUamgszn6I
X211HQiKZpSI/fBJCnWiiDsWx0sLAcdElrta+toHU7oTELVRhN8Al6RHLK1aChKT47QO8xS2SnBA
OMYRblWOt+MtpVznxQJTwnENgxi2+xYM1Lechf1N6od0oYyW6zmT1OsXPznDgHSDFT8MHqnSKdYl
t0haH0fcWCFKL5DOTU+E4yAzNgqDAJj7yrsAc8hHcRYI4uhbV/w8Tn0ot2FbRYyyUxgplBt8ELP8
n7IlmObh7exgEoxlZVvSBZ/LAvs9xh3p23Z79eW+6tqlygP70KJAgekHs9PHFU8SWnhJ/8JF5ZiV
C1T2iW9SNWLtNPV8dfo7IKV4Gs3r1+O4KDtghigdeoLJACl1X2V0PiSN29swOws0a7NPVJo/5CpX
ZbOkSPKb+ZGthq1VMUXNw1wJOAiWwHJQ+gNIRAgVMSiENAWPoKqIQGhJtpHvPmNZlvohQ45QjWw4
02TstZxpzNQ3muUH3q0QNkxArw2U3g8Zdf7+MDg+ABFUC9/FDV/IQYX42J8II3mbm65Y90S/X0Ho
wG3vkURztOZEQd8kPeY31RtI+Yn+BebWN4mFm+jnNRFo7/q/rthzojf54yx3l3YikjZRnKaRV7Hz
CNCFTzl2FGOIOrdIX/E1pYvYbCRI78Uhf6JNr9yZbhwUpecoLbcl/IFCHJq1pvlzv3qPqhQahQ9Z
v5cBSZDtYRujb/+avh1S7ywiuTFJw+KCxc9+Xrfso5rWyr5cgf98KSZM4PfDNkfltcUWXrg/fVzV
2pSKmFgaebMvAxg7uk3Q5ay0YIIB8bcCXfxYyqMiLNIyTpYgWZdFwJtI7eXCX4eQVgP8R+xLaDj4
xATtJSKhhPMY2U6m28rRteqQRXtW28UfZ1Y6eMvB4kx2uP0wQCHeLZnX6Aub+2GO4cocNgGtUhTz
Ml/LTNhdJ2buyIszzBjvgM3ukP8yWilLAHR13Ip8YuFwlOIh37KZ5M7fOrNHriHCDiTSgJtXwHdi
JA7V05owwHoBVO984/Qn1zW605Rc2pqHFwNiodkzlL+4CEFNR81CResuxQIuwU7C3nxdMscEzecQ
xVlHhwBKSBJDwiDjR/yh3bFVAd5hAkSMvAlDQqWkoTOnxvkm9yXb4+lRmlLG+2/2WPySliQu1EHY
wLhd75cXBJ8+SM+uCdG0/DfzyDSCS9GTkn02HkxHvncvV5XYtkISFD6XQJGts5if/gz3mL/Bkvy3
u/vc99dIn6lySCjKTV0fWWte1QdtfJdtHE+RL8G5o5nSvO9pUQeX5Z+C7eYYe3Py6rmwpd2HGot3
HL9t53tambUsnZZzVzvWUCCk5xae3RCx2SAyn/Q85Uf25h9Fh0M5ElorxtTsZQ6HnCVcLoFAaL1g
pLI8DjoGzV0PsRL2fg26/Lq5WM4cDCctWYq4x9a5op2d2JArHH7ZkAp6GCSZM4tKUwtYxc9mDcIf
oLZ2nSCLsOb1lz6cadixeYEKw3NwM6AFNXD0Ubsr5UV8OUTqMYpz0zAIJHrwhiiW6t64fSpw5nDu
bIXVLf1UErIwZxsOJW6fev6oXcg4PzrXJ2Jf0jE5MnjvPYROQxQPQof4n+i996SQrnVXKSJxpTtQ
8O1gHprUoYT2UW47r+s/RKHtvE/sEjh1CcR+wdF4xP8NBZ4tBs+cKfYy9rrlnPRwg99EhH1r+4nU
cl0mKYDk2KjO2hiuq1nYXTKfZcVzlBwzEfDZDAhybqVNtGK7T4KpHgiqZ1zyCbtzFNxqTYGUdTZe
+sJBiUWH2SQx6bpT+sgoaaP7CH84ESMSKowBZtNN3WHFguV20dNCJinXYoC7rzw8evevWuQB5kVp
WkP9r8h9wrtSMzTBQ2E7Tpka4nA/FvxVs5Ycb4PevfqrSOhfh/sgcDqUMTyzNOb+XatpTU0w4M+t
6ta4KVLWJdNPFkcfg+GyMTBKyooHxpsvkrvDZG/ok/asQ2JF+z3PizHTz88Vrn/TDvnWhTnLT+BY
KDox4ovd+iBtTDZr2wXW7iVTi1Hf+SYxwtFGu+NpNohQA04G+kpMvO7CMgZupLZ79qanvAYNEQpq
ORkR0f+YvZ/RZVni0u7iiqIsRnGjRnRr/ez3J5pDtD3E6BLEHPHVNj484hOjPDpdfFI/gm8puplP
0VtLMwNpGMb9l/A+Q/OuFThWAwWrlSrtG7G52ChlpBFYGl05+9M47le0A0ihhbeB9kwHNiybPtEB
dD3Q2ywGJvw/JlKo5+o7G22zywYqG5b5LWRmd5sMfAGnKsb00pRBltRGrvV39ynpdFw4vHK6Z7AU
jwPjx6mKPpfpFXHAyaq2pwLjVXOxKGhP4RYu62sCDkYRgLV3WlAPigkPXaDL2LaSQNclbm+nwbz9
NV90KZ1HMJ8fVmpbcaQSzV34+6pf26KDEZTLZh4JG4SoidG38ZoFb3tfOnh3EHgDqAJmGlQiiB9B
ZUcP6U7OdKq+WLIla5/H3InJcGBXz+P8Kh7vJswn1ZJ6F9alNXq3l2hiBtpBlCcAiRnxyrqkxS9K
g4ek6KOOJtjtbQIjC/PmD6KYuQqCso7LIfmvGI8ReTDJ47vC6ybYkAYGpNYAC//nP6gwguUSva0F
NmwfGn//CLxVWBsfDEq8XqCt+fwVOX/mGFW8J4mzvgNp8f+t4FLC8FXvonPcUqE/9XXKIWPGoIeo
UgTLmXLkBCvYxAOkc8DSr+Y9jw/MJdo0PbJ8PgKBLILECBs28m3hdwrQ0CeQT+z1cZrUHlNsiFQi
NQhGUQMODTnsQnQYU+VRn9OQpzl9zwHyGEo3TSXZgqIJ/edutfRUPegQ94oDhjIPhGNVqFo7SroA
esZFMYPayHGoD6cHrDtTDUhWHyk0EyMIl+92+BIkinwhGH6vRNq+2ZIAUlZhA/CAefRIEIVbZm6s
sWGsdF5P9TME/6+RTtEg1bcZgmKUebWJUts69jaYwWn/IH1c5AHSLdAsTfqBiK/DCnM3bvCI/d9c
n7H8dAVvoPeabgCc6GosO0pyHmpUYp80k5R07pRp32DCwI97HEib+UPdkayZ62FFz0Zdkl0Kr7m1
T6BIF8Qz0k9Nn/1I5zzlF++3/pmI0JTxhmJzy+garjYGnBtVZVdXTRRmNGAG/jAcKceUcc7IhxNI
3fEUKt3qnDFGXvTpr+JgPtw1ze1lvKhcP+P9Xv6KmnugVXlvv0MiBOLXu3/UNT+EMzbtQF/ino07
estSno842aSf3Xs9epcDdGmRXzHJUVmpLYiPFsmcgDlRDdRmwYTDeipIpELQlNrbPMApollpOPWA
5z1XYbror3rS2HOAxoMVXr25xbxsTMONqWCCrLDJAMM313+QCbwcLdGUo60GbD0B/XTZtnBEYRoH
xajsm34FkJzOUmQHgTzdBr1E3vFn3aNNReOKyxfDuwP9syJwDhErq036GHmoYChmt4o95D0ra81A
2l1TdkCUy047YqEDC24M4v9RN0PFC+DIaJLrOa2Rsl/xUL50x1h0H44H7YEe8ziyLFcYUFE8BEl/
Mlz+SKNmSRA/0EPxipPZ6m3hi9j4t14zBEuGX3sK+8tebvFNpoKvig3khbHoSV3JvgxrgaZ2bpOP
e+QOf9NOuHZymWWcxqsD7WW3gK7JRKAhjWGIDPAoz5gq3T0VvBbnFVwFYDgfjOArHz90Od+KXcCF
mgIhAj/fDxmPjjsqkjllbA3JV1xztD8FeD8dIuN+M5KYj+9USPi8uTtmtR5y/wo1hw2EpVh1F8Dq
V6vld3H2J+1DKjIHYaum9GrZ3lHr/Ld7sYTL/kbWoJz8UCSg53PgIrqaKktALeRDip5Y15GHL2AJ
6Cq5V78M5fGa+W3FMZowd/N0wcuHLyBvXbP1PEYDEh50JOm8REdbjCkQdvScLtTsAj9wURDAAFtW
qrrO3gRQyTilfU5ITR/zzShc2UxARdZssgzVDYhCz1/+9e62wB0lCyH+dA6PiPKpKuchIRmJG0pI
yeVgVVtVPaqHUMX/pIwaG2s0LKAPmieal6yoRqy6ZI6kazccxBg2+N0W0l+kyrWY+0c5kE8WOu61
X41Q8rdKHS/TjLjyG7rPISSwPy3O7xvMxiEbio0j03pVXDWh/NN6OKbOJuNB+qNC+UuiU8JvrwYv
XG3avhLZpGCxIPUzeI+6+d6C9T+mAvTA55VRB4L9awZ0y3E2MFXIBrpqesqEC6T95TujRrmD2EuP
4WD1lCp0HSAUOogPujUh4OG3uYOBGJQB8r++/gOztxQ7FsgfnWC7P8YtF2AGM3u9wQumYoxWlUqT
G5NcXay8OtbDL8ivT3Y5eQXZYgFNlzn/QY29+f5pzpSZuUQCijaCnEDfJhapKxTuysyHcjXg/I2Q
a0F1mt6OFSV4jkngbjHYk/6CiJoMqn9OV7R6c60wIvfp68DGukycHcAaj68MC7T4sMKAphv3ToCf
OreC3uPX/GIHmd2l10XV8w0kX3pjmqH0AH5c3b3EXt5ah1HxUfQGgpGJ9EQc0q1b+n4oP63DTA0M
TxAZI0KaF9qCEWL7toU9EAbfg2k0B0wwI2Apsi+LvZ2dT64WHt53u/f+txv2Kjc0LBCOj9rKExqh
Bfm0geAe6d7wNIfalM/t88R4YFKnnGUDrI0swTwHsvEpv6XAvUrFKx9GdPJA+V7ZW/bVcwhzhZIo
y7vH07go3RoYeitReHXAP7cRCa7ry0jgvRYbOJ4SllwZvXl8o8XfZZH12BKrPQlSPwBQHTCWW1y1
4oEtoP5WYcu+EE/eUn3PtQSvfvD/HgvLX+gzj5GH9Y0gMKx0Aro1cronPgD4gRpo0NMqVdmNSTXn
y4VKJd4rq/v6p4txilhW9YM84YrdlxSOt1fUgF+sv6cX7T2+hyEUBzLfviXjMBD7tY3N61qOgpUR
4aPZpgsrps0YxXuYxHn/UoodZ9Ja/jEzs/GdAXVY9s+5gtGiGDak28GCaX/7/5UKtten4nkXq4IO
qyB2InQISGD3Ypg8R7CRfe1y6A0o9Yj3E3tnHyUTpGmeBP1bA076Iv+mX0BJMiVH558Fh3OLmU3q
AcGnLnmqx27B/CkcNJvUT49AD9EYR4H71Mq6qNMuwz8hK+0lFDftDQZ30EP0W822iW4iwtMf+6wK
2ObijfGWEjBeC9D6PDEfuKjSXGvQyuggaDhQwB4k2rd7boVd4YeotoxWYQ0tjKqrErKKEQSYxv3X
U5EjBnh9lt7wDZcri9Eq495kQrDejVBa0g/glJ+Wf9nn2eVLRGuuaPJt0590Hbn6TGlMDXj4dLeV
+e0FKGah0di1Sro8S0JJUoPB4RyXyA/TIg6wOwQMAzBnWbtQxmU+3wl3K1+3tQqR8jdOis6pwu/m
WZSpow5oUubUA2gwygL+o0y52QN+1eT9xW/L584ScSP2dHQTqeLX/NlcHDX51Ch/Zh6jHw3UWvFN
dboiSvzQZ5o5vKDHgaCZ8PfIToWWtpUNBcgljgIswrrU2VgWWfFMfiyyvjFG5MLB/eHibumOGhYN
/Ik53dJq4P0KKrSw+NsqL7zySSrJO+vr2hbWaJgsusbqqM5H95N7HFjtXXYuP7KUs+ESgdxPW3FI
Kft1JffTxm9jksboS30kyoEM+LUXwiZDuVzKAXFWYLSkgQsQY1/Vsh268qZ0OteoTODy0lnSW1uJ
OFHemCvhvWPm3VfGzK1xVnfyiVTeLL+QciKZh4T6z9+8RdTxGdyhiSCZMvyGuIWr26REHb23pj+k
DNtlDH8IV2PZ1akozvDWVmWV/zgMh3h4+ixTqgtJTKuBHzNONjO8lkoj7t845pkijkKLkQRWrqsx
n1ieQF7toMGuKLx0PujxD7xeNyTWgnwv+No8gvyOHzqf6GbAwl3lH9UEBbdax8y1fcqhYTXJGTrD
TBJwOmeZdZ3exukMU/DCIgJxFXhQ3OnJ2S0hIrvjTmGX7ER+Fyjp1Wusa5ahUzHMX6Hg7frVD5g0
8pib8apzYa5xYdEJoek7rlMUg+Lo5L3ig2YAANOXjxrQh7ZuEas1vo3jXnV17swlqgd8c9GWvxar
WWuM+OnQ2uTDiTi7aSQuI5GpV76kL6pcW98E8UWg9V83SBTcEQWQCWdUhZDyYcFfohVGS1MMecXv
+S/aSx6iHpY1xEis7qBmOaePpnwd7sjkbbxTfNy1CdHznBy8S4qEIvQJNsUmK7sYZBhrPe5IbCxs
R6GJoqEWT5hu1xMMKfebBiVmHTYPJ5Z3Mki9RPBr0Wr/IYhhurB3tp3yMe+EUY9L7/EhKaSCAE2a
Hhsy5d89DwFlhPPiQU31LwmftzZM5/+haJ9MjgRCAS9/18H4+Sth3RB9seEOB0VD7Gwp/ZCGMz15
g03baosq/EDrMLccMkTOR1NHH//Cy9/YrM4NFFq2d75ZUAj9vHrV1fSs6ISYCsDkrxcWthdy1sV8
uLi0Dz8LKDTAUWUE6ygRDDH2r4pupWqdXor8NPYlWBITgwmKv2lvttPRSQke3eQEcup6qdXcqucj
gwtm9/j35fpdqPTyekF3+uJNM3OkDSZkI9ngNXb/uSFLX0L9VpqMwapX2sHkPE0OH4iYlgg/HLam
NizABuVrWrLAlq8GHfvW9D+ttAcH44gaipbAAybwK6pvbMpRKltwyPflo4l0lRnHQMTkHYKBOmD+
V4uc3LtUAysiUgJSfOpja+fZa5kI1E4HWhQh4pZs3Ef4WKAnprRnf6SJoQjAvt/kv4FB+IzfecVv
Leu+Q7Fre9VOIxylaL06lkHPoUg22Ydf7cFy5k0M3Vi4Xf7F2Dc/93YEXnXy6IpoPp4l1kIwweP4
GxeguEFxtsXVMhZ7ub25swrjqdwHc0ERb80Z1whmZWNc4VuXlaqJlSaQFEqNpKA0iBbVFp77MReh
rGzZm+IV5C7FGo2PobKD1p+S5FfwaNLTjcWjRJ007DDQ/0zp5EgwC5mbP7OwPon5Lqo+yZrJyi8p
H1IH8VmIfeW7bEM4GSVVTMY5Fd/45gi5+WQ0zL9TIaAx+ebDumrM/F/bHU0ovCoDDqmLXJpHo1MZ
hRV1fXLNmpQfjXVvyJqDbRDP1FDadsguNaxKJkcpk873qmmO7XSQ2v6vHnIhlYQn+IhQumG7MEzh
lg2VeEHzXs6EK/NRPfgV9tVOo74ZMcV7LXYDkRFRMMvjwcBwvmkppeZ9xb+kZdxHqOkqL1ROrtN5
ox+q2FdW2YRIkkC/Oar7usCsgEPFwSyn8sHgFzLfi+uG8gQFfUS9uea/BxQMTl6+/rayG1gmjK+c
lOj6s7jf2yWeaC3tuBPtIaivQe7jqcTbjVSj3Ioqw5yw+yBL6PaRpdSXWtQ2/vVBnQ1jinrwyKWq
N1UUrk3Kva7fDJB2CHvgfQ3eP+1NhyRSbVxdOgm49HYCapkTA+Eq1hQDPJsvc5PTuRTJ320RBWw8
17VUjCItvAyhertEN586KQErdtyGFaVVR7J19WmDANuNsrYHEiUKj4eb0007dUQC3EhJOeZ5baDp
JCoQmk+dVRPzC+ePt6wP3QeoZduVRSc4ILecw3DkzR9lDyjB0hLJS6iSXBblkBJg+Z/yu+EB7dd6
4WO0V7CodbXjhwIxcNULcuCL4StNwmDq/EDgD98QPVAvxzUqHOza/C6keVknITru6+bLs/1jDg/L
bYcPDgrQjrrSEsl5VkXjdDpFkuxtWbrMT1JAAvTOXvsDNNoTpZteLb1Qi+90IcpQK3fE/luGZDnw
omHhdKixqvA4S5xYPIy0mrcOzH7i6DBY7xzrznZ6rqVEXr3QamyHDr7juV6aYCONJVAY+ol4wZOb
teiqk0WRdYlds1S+458WqgAnZXJ3BgmoJ3hxx+j8zaGNAcN5OW7tImcLRQ44J6QvUMi3eE0Pi8ci
nsYa9rZvWpwKMTp7yOfQMl2tfeLUgTpAcYrp8lBE9rAwEO/MRm15e6pfFcQnEeVdrvQGzmrm9P2t
MNlFYuEPwb3lNrECh9JmNuzAJQr2bk2o9Zs8I42mXdexXKptnHp1iWy29V5/nOunnexQgM//hA2a
JrN4HlgCyfkHBmU2KkP8VU5ZbffxptZLH8v/AgDmrVCfxtCxKqyCm+lClOIbR+8o5tB9FIsvqp3K
Nu1XFCPa0Lk65Ez73hA/mElNlG4qF3K9GXcV7iZ1ePbhbNaG+AKwoPZ2PvzXNIXTA7YSujoAC7jn
TH0LPjKs7L9GQWsuD17OUUPmEdLgJAMY8X0UltqJD4erjAn6Nd1xQzd/fd8zYh0sZYBX7W0aueXN
HfwQ5zAn77xKxqsQIqsMTxfG3QaO8QEKDL3j2vwjSe9ZFm+swUzNroHXrOzS92wwh00/Zz7W3qxq
ZnjgumKRnReAMCnkWkJ2HngWHanY4a0kOc3hGa4GlgPyk9dDvNUpfUePoTVZUNQ9NfPkiVL1yfX4
PmqVVbuLxGORYMtPfXAQfmXEYhouS3EmncyILZHw1jcsrp/j8++/Kakhovjt9f6dPFBuM7EouKXW
6i4NmP6NWInvgYz9thbk+E2RWuvLrqjIgivT27IaeX6zK4kkpamK3hTN3vdVZGoKiwse7IbXsT4j
JHM7eIxl+eRxcNTIs8aueITUEiQjHn89BQxZp5QGGtSAeGuLOGCTm6V/Djn5Xrci7PHcFE7VP9Tx
0Ub2EH9e38PO6wZl9HngRQWWGcxZXHHyUEaaFBfAThKMW8xZKspUGMqbcv1NVrEk5TMGKX/dfKZm
9/7Po9jCjU+al1fE0GIecpUmht07ni1iLoXpTRSK+YFcQWBaAliQFcelosROjrtIu/kHzvIK215C
Q7CxjDSEHeEcT95V3/bmO07srRzBANBn8oImUqvkJfjgoy92xSRmF1AZ9Yg6PDz/VA+/pTL+I9Vo
3vLBFSI3ZOxRYYAVC9JJRoOvZ4G5XZ8uEdIoU9mnj63WvnsE1n0Ixt3Pr1kshUW0sGkLIMkeVVAK
4hs0OkJD4Jowc6AjO9UOH0jpmwK+Bt57XaaksGVQsG5OdZx9+jgdKFKxxdRWC/DBTESYO7Nw20mQ
eh6C+LOJyDeD6L3xqmOGADtbkkQCO/gV6+J7yLn84o1UPQhJ1ldAZqFFPyP1amUpUZo3Dwrk2Jny
GLEYZ3LJvpxu5yP87gcbfrUBwB9sd9bCj1PsPN1cjau9p6DuNJgZ+N4ui3gMFwpFsMsGmhcY3cyl
gpdfmdcw23hG4yOMUQQS7vAH/lr7VcgWPmsQFaOlueFUJ7GKv+kxEplmPk33/9axjB15u7VSPuOd
Au2WnES0xuQRTaSNTHVZG1HRPpHRxb6evbYTO+UmJ9893AnBW8v3HldW6e78cMrK4jsw3DRc2nnX
b7Cfh0FsMD4z+R3rb+6yYGI7El8XcUKKrnE/ymIGryMXi3MXbZH13UjHuK2ihmzdWv5daf3resGu
dkq9SVQUK5jrMJ8+Bt8Jt/oNYaGOVhUmfGAeZO4Pu9BX44sewox0S6/L9wzpWpkGvBDupXFHgCXG
axPRD7xkFNnzg8D0oaivsB1Da6Z6VRffyOUrbv3h9bcpZFLGZicDVygJuVZpsi+XHCEN4utdufyZ
b12D+WEoijmRBiKw2kvW/ZonrwraCJGgMCnVxry4avbmY5AFbksXS1TxUUa7stDCUiDLxv4EthxL
VhGW/A7MVSswgNgTVZvtjZPaj3jvo7vQlrKBkHmK81DhyIF1m6C28LHAFuM3way6J3hSSaj9r9no
1EiIlyCYXDor4N5WIs2fcXEkY7VsSPC4DlpytRWA74qBtXKHq0VnUskG14BHaXjnHsbNw5TmqHGL
2fWbHf+0m8vVuzO3KDzhLyiX0Cotj8UscIyt7dw4ICaT2fWiPBqoGgzlfFxVNmqdyJj7hXZ1K8me
epF9p5dz4BtNJbs3BblR/wyx/XeBa2PbPHG8gnbSCmi7RCsPD3tWs74lgjTHdg6XiwLDoSRpYldA
4yo86XPXHKpCwWHWOrv9fsGjuLAvCh/sOmzy/arJHlhAQeDZxjLPIhFzXv7dyaLLn0QjMeJSf5dR
gn3I5/7MNfj9m6rDo4Z+29bSRhNtMgKQp3eLHrrD+Mg9ObHHJB2FUt5Xufg7JVjsLP4xdOyWLuye
+TgoI7pSFl32jLubg6xul94yZG8qwrtHDc9CKkomKbKW5CJMr4XCVgrJxlVT4pdja6YfxdJav360
+kTLJ9t9FLsGeXBuEOAc6PLeTfA/GBWs3GGKHLyI640qiwJkagLuWc9MylnmqR4obh5uxTu9idXW
0UDQQBu/A00XCiM0IKmcTOVymgZpwxQVgLyKOPKoYYiUFmBYrQo5yX85u7QkEeKEyWkNYgexMksv
YOCTWNjoz7z5uecKG9LKXBkP4TOaZlcAVIOo/BBwuKAIR2gfaptu39TyQTLGOo6lkekG1gleSIJy
Km5Og4/AT3dkO3mp/KeeldCqhiodq5RXYb7rvp61oZmHXM1g288SEBFNNWq4vwC1eT7k4Dmo6OoZ
A8wpzaukoZocHgCXWkk/D40KLOwk/fRkIMYPRzpIrr0dMH1iZondeVUWYyvKPeYGzjj7GkcygLJx
DXCoQ/rlzJnT1yeKd1lZYL0+/ALOerOCL63mXeWvAiBq3c+tte4WjaNuRCC6/XNgONJhiVNnemxc
kYi9lbw73Ewh6WSR4qO9IkSI5Tj1o1EDeeVKZGGlJAUx1jvAxHL1vAU5HgoEaOuTnabBzxWiS8Sd
ASGQB+bzxecoFxUqxo9qYHW6cFh2v5+KCzvkvF44jiy5GZ+CLx0mir4B5JmwvS3/zuIVhmiyxn9/
PbAZJArq58PbARvhcTQhb7m0EdGPYEwJbleKKcZKHrGuTstgjUt2gc6ge6U8T3kkRTpeZgveFDRl
4enRJNHjlv+LjyRozrKrN3E2nSijAhXhYh/hci7r9UjkCLszrJY2Xq5b95doxoZVAPBkY9emMfOr
Agq4Dn1wPDndc4YQA9XwFsTb4mJTwrFXkdrD4c4kv6z3rCN39BVoLpdfhiDAfQ0phomewRmSldf0
tBJQu6PiE3yaWc5POoBCBEwaYlNGcy+TVjcCcMKKx92o9CNnzZ6hh74u8T5CxaG3MoqdUZgqJM1y
uSqsHtmaPxgkxPuxiWqNVP69lo4GNts8xIxqFjDDTJVOwpywgKOPApFaRXGTEQ1lEY1zV0UXkHi4
IJobVASAM7FjadhxrLI1VrgGL6n7YhSEenn/3K1/vNyGqCAGN06sgMHNmlHlXkI123Q1RKB5jDp4
osVpdjtKWRewXueyQEqHMIn17KMeTS8q77Jj1PyhFctzsgLveoQBSESwvsttjXPD/VEeG2S64gtV
xb9Vz/GXPUGstPCmn6huRcM+XpqHCnzGwMEC/zkIwJDLtSt1VvC28cFimcre+qpigsKy8nwXzvCr
n0GgzeB5dgGSl077dtywhLbED0Jyrsf8zx0hfnfLJKUVPeJZIRRuBkyjcPFdMsI+jeZExBlxAqkg
AOhBjjkUPVJOT4ZvfYumcMQBZsgAsn9maWi1CqK5vgd/MVmdFctWFhm2H/UIBWZdNlNaSMKHY/Xt
U4WhTufG+Yf9B3ddupajufwqeM085P57iRBnb/phxpBuiY9aAxAUC5aRytp5a8vwln4GnaYgpus2
yMEiRPB9PjRB5HMlKrUpm/z14XmH1SM16krPaLgDMgu//3A4UrA3DINefe2JA0sgHMRBl0rGyRY4
NyA0FrO97ai/vhDnNgO+ad6yV8xAUlRWDbrGNnH+rFk9GqRuvw6HvRMcApIXNrHwgPMkcCAOFSa+
IB+Whx7ZOaaVaz5sRwZfp/p4Zl02u3gyWPEGDo+qjaHUTP7Xs4zS0xzIpitTRTQvCmCwb2fUH7Hf
mY5qIFdKvUsm8I4VGXIDzoNfksqFVZnE00d3W5hI/B0TItQ/qEiyOQf5W7oIpOWJESJD8Yne/2Ws
bOXYrKcUoAOQPVaZTbbULZH9Yv2bS2QkYTZn0q+gHlz3q2ZYM7bcHu2e0sPbiviCyPFuBqo4Uc5y
pdlF/0DzdI5Pt90R4yVd2nbeg0/B5Vol/VwariWMT67HWJ5ihMPVQG4K/7y+0rr43Or/vJOmXxQ7
LOySFl/L4/iJW/WbEhyPolGVGuyFJaTSiAwQyCWtd7CzxhX8SxvSFIn2UQDtOgHiO+nQ+Mk0htxU
pYRe7VCx6yk22P9b+cyfDuq4w7T5PVeDO87h2togsPJUCek3O3/78FozgD7FWwaLinT/pd1gV+ik
uVit9aSptp5Ka8mE8+DlU5kwqV6tMKLjypigPc0KTmeK9GVmgVVE0LqWYj2Sw68i6uUSn7tmH/r8
9pZpfGPaoXJRsvaohplNnFjylcjuFjd/rkYtfxd8sQn8+ZUvNhui6Zsx0Y+NRGglKmS/Q87WhRXL
J5GpSYjMbvC4VvCmVUPjy9wijaNt8I0ECTuJfI88nkYVO0nh4Wnw8marmXI9Gjmp3mfO3HyAUjDh
wqZsK+nzHhu234JskuPTOis0HrmvBw5uMbfjwuAigL/DPgbuaokJqIZ0ZzDs08Eui60j/e2PrDmA
M9jNpA2mHDMK6x7N+ar8/kip8Xe3Dzeib4YXFcyhjmi0eureaVxyTQTqE6QBmtUCm/utNqi65SYy
tPntHzv7/3Lhk2ANbxqCgEmRl3LRo1KcEAMtpzBJRV78rFo86a7NgJJIP0io8k6xRoUgRHeOcMvA
Eg9QUaA2PWojj6H9QXKwflwNZSrlT3LpPGFGLAK2rl8u2HRiEx0DPJPgq1+tnzZjcT+zA/LY8rW1
TkO0ct5V3dtJMbcRcyRzVjefO93dJ6Sc9ZyjzF3jOMqeqA3qAwB5EWGUyCQuucGKQeGVXKHkaEad
+YptSqq7FBx8rUscC/bRiyMkqPsDJ0omj4R2GQdGpo7DaY3KeFvCc7VcIPRUtkr4zgy2EAiUfDxu
jZ+AT9S1VNLy17W5wyxuC6n8N7MZHfLpQBfEXjsnOxv10EDNhKdYJz6ddgoErtu2G74c8RWcaaZ+
AyM7rVpV8CdbcEiZCL9nRkfe3BKgIdpA4AWGSTBX1sHANuDwvZvWaEwurPR+QQaS8qQkJb4DIU2O
1dOsBd3xp8tBosN/vh48upD8Tyc8ADq28k2ahMNmWvhV7qteF+QkBp0E68Puqtd+bLSyl1nCq6C9
fhV9ChPYDVhIQXHeCc/XKU0biMwUn8OslYLmvFja6FnXtgU6iAM9oHFYgBt+mcXJONrq3AOFAYpM
dT7y7n/1jIFK78YwJ4mQT1iYgf5JkXWQzqmz+jP3u6H5ClTX5VNPCanfEpqQzq7rhsBZG3H8043N
8P3+QKB+qSfVn3LwLth3kE8qOaoGvutxpu9Y0yPWVvfDJIJi4RcJLrlLvSNqUoui52HHOCWIdFFJ
YWVA5Rhr9fmtzw2jEFv2wSbTdPfmUW7D3q5jXsfP3Sklzb620RtkBPXpZWP8hzOGYdt2DrPZuI/m
GjJBvkswjZpZ7ksLEPBLjZt1O0tISDjcYCe/Da7TwZqE9T542vi97MZ0tf4+r7KulCA0dJ4NZgpY
Jx+J+SEmgMJ36uwa8xoNqkCOzVzTGF18xQNGoWjMZzydQyy8UIwyXiGjH47pyBVAKscpFIY3LYZ8
WPz3Xyo+zI+h64+d0IDYY+en4emPWfhOJkF1xWO8RnwPX/zD6eLIv0CbiE2kgqUZaqhyZKwIZ+fp
3hFOK9jbcpQuPDXhxkOCsevvl5D7hUy8cBpMwiIHyuUgTq1jJPGftMoCxF5VkrAYKlWtuksANsmt
7gDOnzRqX98zXe7vJ24TLKNoqMjeREMIiT7mpCSi/eB7x0S9tg8u44nRu/iDuI6OUU0jwX8CTsZA
ovvraeXdhgjjR2IWIouqrsjSnpkwsTrKpvMQp0SwL1m5k1mII9BEsbwoanProh2Ns1bQpg6TY30y
kXTj34K26TpaNw3D3JDEB8xjUrotkTV2/zBwOW6mmdLDCpHZ7DVtSJF6XlIHBX6ueSy3u5G2L25r
n/VUxX9O5OXj9NJ7hzHSphKot9CkjqamFws9prG9ooNJjV/VeE/PxxHhbZZIEOA+NL/CdjNyZMYn
ox49MWmy4c3bO21uu9g3QJdJEnONWj+qrkiFAoDl9TDGUdfJCeJbivEfa09/wt8tD57MC7i49lKG
PoBCsRVoU2sgvJ069AJc2+hyiNl6w3GUDJ8vP7OiD3U6xHbfRa5wi0MnZCr2UWni3nhYmp4aPmjY
L581f3goiLD6xXaRt3AhESgXdByav0IZXgCXydv9pfT9/nNXydfdga5uZO2dj2vKXKW88Rww9shx
3Iqy6nb60cEP/WOjLzm0dhGxMPHWwyjQV1wWapcCjKUPKnwDmnSLdZlVlNVVrPOMfA4izQJ4Ducc
w1sb09Cm5KXxKZ5wzFUuyB2Mbjj1DD5eEVWrMGkx+jBdhVyfyNR9Lawmo3hsaND8+jBJEdusx/aC
ySUjM1v4S3OpPOB3D8Vt02TW0D/H8M9Xxy+s3vxFbfl3ro3KQtqr2TNiiC+rT0Aety5ckzHJXj16
8vOxWjUXAM3J6fqSlfCpREk9GDFaQoj/dH7ts5Vgc6xvMgCNQZWzDXULgx6TUV94rHObcWaL2Esh
avKC7dlARAD0eJ5Q8VdN3Y+5QGbcU4CZZjx/R7euRbfPnP4/7n91uLlpKbocf7vMd8f1MOkFaZXe
Ak9BxOq6HgUOn4iG4aMTTtNK6D56+jr2euLMLJTlbE/h4mG81pfmUIvLonR4hgBueQifiV6gh1gt
3pDW9ukWSLhRjAzOmspIxUgcpkWOXyeigdzhUyUHlIOS6QThrTprs6HsP9AEl60V616Otezk1v+S
3oZ+DchmqTc4LIM3pQpEEZixQ+bKtw/Wq605DGBVOf2XX0pwMgRsN6YJzoDhMdPwmGPc5FG6geH5
OpWOy8rt64Xcq9Uptoo+B//pTOWPNnxSe0TP/tbf463rSgHTWT6K0At80tVX4FhiSokxFEmLR4yO
IAA9F/evV+vZx2oinsN7Tex9cX/MQFtsJPyvJtBUTCHgqwiv4dhz7srnnXS1Be9iDiG1ZuNw/bhr
YBIYGw9p74IOwLwE63WhmVTN/Lpqjc8uGvnagf9GxG1VJx+hJ0Eb2XXTcZPZv1ulxja+JwZHiUSf
zIdJ5NFcNcYhf4IHGWwaluk9froRKEthG96edi4gkFgXiUfJssOaIRmyq6x/haaElvV1HCHV/AAh
DHLte5TxkmmDOYHtQOvDYeIvDV30RQ7t/dpOQFWD+es4M7ZYSTf8qWEhcqgnC9EQWBcPcz8r2JZS
a7TgvcbgHih7BxsNKUKw48RLUkzNkzagF9Jx8ZbxLfK+vVQXNIbW0W75diRGe5w3/nZEVPjExlea
Ctq+AVMrYerzrlR2EEHSYw0eUbzO+v0T/Nrgz0s/tqkEeMPbr/fO29WdK9PDpZh+te3USxWwFtdF
Mw/bB32PTzgAsmRLKOgAfnwTnsO3xcLwQH/sNCbD5mxW4UypeV7dnZVlQi1ykNZsITKofb2mMTsl
Gz8ZDw9i3i2atjLDyvtQaR8lfpeRKFNu6HoS0KpgYt8L75bSgcCKFpOfrr7D7BWNscAiXhZxFny+
Gyvo410Zp9RJOXmXMVDtn4tT2qIOO7lzjFU2PAFp/9Veq9FwnQ6D+gpjjtcq7FVGprwdCkQoiO+D
Nmntdddu9jTTwnBjQJwfEpxTUwWJEe3DcMU6/H5g9AbrJgfp/dEZQkBl5kUlPkwQnLLHyW4ymtza
tBaxbZd+Q+SlezW4hQnc1tPQCcOJ67PEE/TkItdfDoizwdc3xgw/kVFJM6DMEDUH/+wLziXUG2B6
/NftXCdPvTEt3ulUAhFV3DYCZPDEywUyhj6a+u6+tjcjoUnEAz20klesegoisc5EpXTs5MrwtW5C
imhehc6fbERbXcB9FfRu97DuMiptaA==
`pragma protect end_protected
