// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
bG3ub11v1ry5LCcs8s+rhWppm6x6BNlJd1Tg0m4p+MK3Oydt8ufuBGIvdE1uJA5drIxVVag2KRqS
sRfjGs1lnrGFE+4Mpnmmhtlm1CTWhl4dZq4qSstimGgWLl5IVVut6RD2JEoI5tw9pZeXJTP+Yoy+
5hHYRm6UUXoEnQCb89nTtaDWHE+nW3MPGlxHpNfru5BFrC+6gn/iFyCJnu8gYB5TWspiO0KLe8D4
9JvxnTeb8bUvYNlOWExG9F9tVZDrms3g1VZBYJ7x8Coppnne6KD9lZMI+8ZNZBC9XnPdmmZHaHfr
SIEFGplNlQBNPjfeSOUpSmP1MAT3No3Dc+Nz2A==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
zQ/rzC1g5R4gLowFKDtR7gc4WKDBxbhASqG/X4VlEG0VixNMbXv1c6IYK0XOjHQ4WF9iXdLhyoyf
9f4OGOkqnFf/ywJwA1xEDW9XQ3ko6HkmxKNl9bqIzRvNKe7b0cw6WS9ITupCvprtm7LACrA7tUaa
edCELeUHOdZQO6BXlE1iNgPNvFjSqeYVGFDsqRt7oy2J/k93VpRXo5xEkxkSEqeayJhqjGsrEIAA
3qtXQ6wBya5gjwGRGCIMzscsoHtVFylQkF2u+mdb0lRqGAM+15bM1hy/fWhSBS/4hKJubhZo2eXi
Byovg4NVF6Exel5F0VfGRfugFo4Ssx+Ar4tf5f6tGoWtp0U6XmdAS9qPrl1WEtycR67mzlag9J/G
fDp8dLgf5W7OfDTD7rnevA6tJNbOV2i8WoaoxrxxwIa279Q1ZwvDyQX+fZUtYgTpkz953ApxK/b6
JTJOnMq0titGgRqhZdcRDcjttxlZn9tEBer+7ODXsTOpiRzWRmrlgV2hSuUSuu8lVgcHDZ3fB1Op
zVU5vzZk4a2eyHYDXWDbXLmLcw2RHodU51rSBpBNhKorndv7g/59IkP/YjEr41jicQm9h3ViBMlm
VA0MDc7wd6LDsi8dY+qlPaO0MvPZqnAs58kUg/mZEp1Z/4KHl3TwcbsCsijf8FJPs+nU2fBJ5sYu
9kaJWIaVGNrc+6R8bQiFnWeVYRH5by+D2SWa/EKICPF5ry/gjyQPs36lqd5lT+iPeig1nG8z5cyT
XVoPRKIT54ZCOZCIXT0u2cYyrgwvH3fErWY3PZ/6Y8/dnmvmUGnCGlrLpCM2jEOyCoxUvLVhYJ4D
toKeyMwhWBUBZR343qEE/YisHI3Al3s/c1lW/kLNdMLLvQdaSQUkvlSzbHHsz7BAaByDgjAgF+lN
GlKVrjngzsqzPwapIRIUmOcIi59ku85Gy382Wwvs0h+duriMVG0tbMfuVZ5COo8mFpNBA+Uj5S8d
FFGKo8+AB40i2PcMkne+UL4h1+DgBJkG3I4UsD6helaJb5FCnwU14daJlLmjN8XjHyCv9B6VAnul
YNkBpPFGIdt/3yifmpHcc+k4TSa0myua50dv6fr2kE1e7V+adKzwnewJqV11sItdltsS+ZONgD8r
SHu8z/bn1x+2ApNZ5WgZrtEOjL8rIXY/WnuR2srt2dyadnHezKIEe8xvBBzlcDotU2Fjz4MyFfFA
l9MSnlKTu7AtShudRi4/sE3bsKVejjjblDnBUTfbdPYpCsZ4arskzRlTqhLBbPw6gjo9FWGiW4Um
WN1U81n37lgiRfEYBg3nRySnQY+eZNhtpwjtTRZDEGFQzhTWndSBC0lhM+AV0XNTouqee30P0C/f
WaajpzL9uiYUPDpF4/LP743HBePla0bNARIQ++MKe7/Y92sh/Z4rbbl+Rco5YHj4l0upimFzIF//
ddqfUZ9xG+zbe7HszLZuWGnAT0ekWJLA+G/CeilFi2u9ml7IJeHLGvDqVAD8bty5TzNVIbqL6lJk
LEfz0QnD5aSXInsDFVZm4B4fqa7YIkW/NVmOZLBtMR+boxVQoK5GbjFNfCvXXGVmikeOc3hVhKCE
n0gXK0s8MubSeMjVvz3tdROjZNFCKM4IavbKIWCa+gmEjUQXD2RqgfP6ODtGrsFInPpIAXJSSfTn
cc5ca14nfg59cDdfmBCmZQ1xTXeDOK18Akn+Oylmn4b3EH/h8MiIlNA/jU2KsZA27GO0dGBPKYjN
v0H5ObpTEHX9VGoREkKFvbw5sXBNLN3Z3BdlnaKHq9ZBkaJMrULk+PUrpF0X44TNe0Q8+1UdPBqj
lkBLMLd9cD42hhh8BmTuLL/r4gwjGKRjhySUWSpPgpl/LvzpZGj0cbcNq9dYw7YC2Q3hdzRArs+r
fQARfgnx9WQzhx5p9RzsP5anGIdMAyOOvMBQY0V+E1s0xv3k7Ozp4Mzw50OI+0SQv8ZLEmY0tUos
b+M4r856Q6iZTXnx4QpKVcKS47HORmoUFdFF8YT6dZFK8IjGE/LhWVD1qbELAvmPpyPeZ/V1QZt+
EL+rzvLBJuWvHrPYBJL7NVgRNgpVkPrT5uYOf+BVqtpClSQ2fIAFsDLcv0uJvcsgmOg+AyC0+8IK
48X9o1Ey6a1OAoQDphwMUVSE24ncsegOiUBuCEsE93Torob7s9hlBS1SbFwqizb7wzB0YG8Rxa6F
LquO5ge5nKIuCOZgcdYJHHSNF4ti6+MZL6JLYHzgX6jeCyw/omMkYKB3CoHggYsk9xKnuBve39QE
yzpwrwFuXCKn7m8EXWtSHTKmC3bufLOOkJItUaxTxuQ6xqeaE3b0vIbv335Af6EWhWp4/gNICd0h
F3598HWhEmfIG6mPwxAYcrZdPD4FIQ4GDPF0/7J4u/RNCpqbr9pbQDT/JiAH4RNf8qAdBQ2WikRq
fekcIuVqrIjnDTlHIuXEgAv/tbEbY33sc0gHwokEMyH+VL0MIPL5bOpjZcGo0DIWoZ7L3h+4WAnZ
ciQ5+7hMkKTRsDZgKvPhHshLFvhyaLLvXIAN4PkzblBTnk5hOgoLAn6b/38GgEMsgE7vrf5Uy/Uh
gWGobujvAq61m9IRZlRkGRJISCSX07ik6RUQZYQ/rfBUDJDc4QLwbID2Suz4eccxVlyyHweoIUad
uSj+cukbT2ZpM0dF1m2l9Mb0KgEhdpZh7nzJ7MsSpZ1LF5tAYRLchqQ8AO4Qas/VyYpqnEJWBUhA
OFrPBxHi25zWeKzs9kb37i62xQbWYmgETnfYzhVkcqX1xdU0h8xWjlDRTbPcxfeBNBqFJkMh95+A
mkTlLRVDva4E+DGSZBaScCV0FD5XgP/fsgHJ8w+19mfzygQt9mZdpEghttdlyG+nq5jrdrwVqsn5
SSMKV57+BpfGdlFoAbO3lItorqvfb93PiTTGRePxOljNWg5J4BCs1WbK5RlqtQYRHxgQx4DdrAJb
kAyFa31InRjBAz57eig4vAw1VcdTs813sA+tM86IjAZzMmROYmS7IC6E9U5StJ9GvGvbfkBhiL6S
Ffnl838sKjockVH7+K+XBsWhkLxR5f5GmziOxtzXy3uk23xxpPAnOI7OxXn/gLp3+qjl/UU/YtVE
Rc57QBpVAOwTGzjFhP3KtWUAoXoyEoy86WP2ahAIXrLYVwR+X55DGpCErprEClSF0emyNjCyl3cU
6e+TR6aRbHj3vZbjnwFL7xBlXl5HNB6I8apoRFlZIYvJXdkR8X3QgR1SURBPkwaXn6DgrFGZVFzr
v7fdq5+1hK047wSZs9hGnpf/6unS6v+oaavbrXA02JS/EcBYg1UmWB6ppsdYJGgzC98GJKjblq0v
Lv6YHsGChx7wqLE9ftyTprlU3mu8p8aC8D8ZmPSsQL++MqYyzbsMxKXKg/A82rGmldM8daT6sm7q
hUCa0syc6NzES1Ycxk/dRhp59wG7aKhwLzGWYbrN7GLQLAkFQcNIRDsn13CXMdOqrXd7CVvmXy3y
ViSvO/3QAO0hA/SLkB8XU9rjjLBpbq/x1OrYufmDNAkPqL8VLlwdgi+9DWVkz/mYdsb2uwhKJjg0
CEOXlzOX/maiqKhS8l7k3nafPuSKxBHv3faTA/dYW0w/1ZZ77iuMGp9PFQ9L0Paq7kP/GAZUDN41
T/lnyVyeXN+CcoKqf6l30FVteUJASlGdgAgXzuHMGBOk3ZOUWjckgvF8mcHcLbLXz02jhC018WFz
nrb8IsiLUjAy5C2704Gh10Q1LlloBFVuoR+Tq+JHCu5RR8EK5jwS1vXDBATZ0RgkJ1wOBM09WqcJ
RiU7k0k40tWgk9b0zF2xDK31jcL5tiFxSQBKDffu6NPcEn8Rz91gpvgclnK9hhx8e2KQ3ZcD3tVN
BAJbHjc+4rt5OI5+4/Xl17FSB/Q+b3kriqYbcwzmPRjT3LeMsSivA9GXuAV5umQHNenvRd7UdATL
e+LsM05hGLhIskmRsCLcCFitSV+wHc//aU88/QhpYsS8tTir7I81D6xF26fgPIElv8ztxBpQn1S+
sPJV21PusNx4w5KsBT+V/8wNNyEYZ671uG8tNzpex2VmcbPs+xOalJDn7EK2Bc13ygI0mggU/6HL
JrIwVmFwWpDKDWZ4BXrUvALTB4af2n0Ngj7flBMXTDjSbStZYuokT9GVEkC/h8iYKi8M0XJ+XgGU
AVB8rPZTNZxBwgzBLRnsNuOhETcot3W7DonPGyTicPm7k2w0tOGm/57Uql2CPExeTOmErOiQWK4D
EVByjKU2vB8pAQwLz7r9Z0akteWxirSX9YkSH42nwsbM9n0ZN6xtRdNx9lrMFRMMWs263lDFSo/I
+wdem+dGDv/xnFMx9RwwhfEYi+nU/xb8vbCdr7vwE9Ei09ICAjrKyqCXoFhE1hrdOUUvZpPEaY3x
xWrqNeS7cXhbjfihpRi95q1Ga1RORKLRIiZjaZVs6q9KUtx3B4NVCs4LwpWl1N6SrxD9MQuwEdMB
cC72eNFBtREeq6SPOBik1Lg6tmMXQpjw/KJppWqqsSclWCOMr2NjLaiTq4ZhYqSPGjOdMn4p7gAn
gWF9/ZVzM4aHeE/KF81LNw/awKIYJKkNfYjWqIg81Lg3xoKO4dm+348+lFYntWRV7bZ9HGtMweXa
yNS00hIBQ/Yz6tt4a9XshN18/CuZZkypGUIzwTGarwCjkH83VgGeCvavVp7Kv9ZYlmIYOIW9X0I8
8I4HIeNJf0jjN9byIBgYz/E2AQzBPvPDYSmzHdU1X3LyGB7n1ghmdKFO/nZn/NiNfn8h+Nuimc0V
Psy5ziVtk9g+QMNaQ1694HaFqcFqZUs2n8mWM4l4oz9NoCgfrt9yutiMU7hIOTX/piYD/jnF0zRg
ADXMVxh+OzEbdCq02hdPOh8AZNnjb92rrIe2sifw5qOdOhuKeU4yX8nw6LUqoU4v6LclJO+QzrEc
SyiF65XTYpd+x0t4cfemEbEzUeaoenn4Q5S2q8wB184zaTKDEbzvNvf8vYdBHUMQVsJZZQErex1f
Cimmc5x5ZVj0rUzrLo2LuTN0kcRjkhN661SJERplT5GwpNF2rhP3vhXkXFzjey8woX4pXiRFYFS6
Nhnetond10dN16iA7Od3AkpvTZyevnUqHcRmFEww0wQzRjMVS8FWXdj3t8WlH9twg0OvFYxGn66Y
KfRAOJs3b0KUZiZm0yVIbaDoqzBqybrhudwlCpntuk0OvvCbq51i/5m5EBmXD9Nx+q92UrzOBspO
4zxwlu449wRNkGR6yOx32i7ArTAE9hh35Oufq1d+na+cZd97vf8678JGgmZOGsfc3Vrc4yW7Llah
M2+O79ODff8rXSiaqnHMaXytBkG4bV4lGyuFTizGEOwddoKfyyefMGq6WIAZchTGEtMU00+VOIJM
JeHCK67nE80LxJntjHPB2dtcj6N4PnJ2fo+ah465AY48+tA8Augbgt3bpMlqI7bnO+5NZjEIk4tM
rsP+VkUBJhpRv6QQVWAVjSUc88W7JzKqe1rOzNXIGNuE77xHnCEIMjGcOTHZEkt0nAKxFfqlxcu+
CAB4pSdFB4mKoC0TVBWfMWOf6XEGeTw96YpXHWfPYSP/gfWbjdj1tw+CxA0iih1qmnJmuSStqaMK
bjfGNaViio4jMTM7landf3bQypILcVXSeEd/z8vCm+yJQucCUYn0yWp8EnrdyF7mO5w7mFqWbbfI
y+cwwVORK8yJ1CrlgNGRh1lMsdRIOgvtioquw7mdF/6egQv8HNdueuBN6RiDbk7bytOVq9vxLOOD
o0Dp1KZo3WuPAfUFJqSKv6Kjna134OGw65gu5A9Eb78szaZAUf7yBDu97196yX5vnSy/75YTK5gI
FkTX+rOG1FemmgdZ1V1/vGOME0h66mFZO6Zo713oHT7gtPezmGE45ekSjR7MEZNjdveAn8sy5YlE
lODv1N1RN2dkf+/ZU/2yFI0zudXNgxCJ0+8tWZQHpxgIoMzNwDS6xv3RjbPHBEWQGuQFBz4IXEna
0LYFed74Ad3KaVkBvJaWMNRG/PXhP744XrehOjGERejaOnHWDnNTzmIJtZBbhLDLarfp4fd6fLhZ
GmZ+calUWDB7RdrXYedqbZMemC/SsbE1s94qP6+VZpsp9U5PzW5EnzsZM4p8vvPHJwcRBpk3cHYM
M5W5azAG2Xcp7UZdsRTYFDOG3RoZNy0chleEIhYMoRovP/yUVBdTmuhHko323Gn1fyKdWDeX1yS9
kvPuBJ1LH5OcnN4Qbu57/DD1B9oH2GL1DkHkekYTx8GW/Lqfo0HUHxvAirEvyehmkcnC9E6nrK5F
ktPVJsB5EDOcKoBoU2+QdcZcuyk+Jfjt/YMkwbCTC2ZUgax6/h9HctZtsAup4vP/OzhC/tWLsL7A
qdavYhRhpuBj104mgO4hfX+wp877FyrGyoYj2b0Sgpilm6rk43QLk3vsLspFoywHYyCYDPXfbsuS
kh4Wiqnw2LYboA4csWJG65VGsNqaU85U7lJUq65ZN98nlj1+ptRCf0EiSgf5EjtM4guGTxk1H0/6
C75MzIMBapygcuciYF5XCjjicYGrvCWMJs1+mHchM1cC6y0S1Z0Q4cMbRchj0lzESeFFjQ77IfPz
/sKwBmrqsWwSuj35ACBlan2mHJRqVcZtuIva2bViOxJWXTqyMlOkgiLQSQy9Dt/siLUWfqdb3vQI
MD79so4O6KnS46jhGY5zqqz8qnzo/FhyfmjwisfRAikiD03DsIe/c4+M9cfuSh5Stqjb62XU0GAj
MduIOrsdP59BoiLdKm0BB0jk3k3Q2Bdy4XpCGwSvcYfLYkMGjWRZHm0tutNOFo+w3zeNsuiwmpNI
BwTRYlJ05SGl6JHo12q4DQKaEHK/0ODO4Kub1Kv4H4DQCYdkGQeDAQnpt9FXjBay9Ozd76NcMWej
vT/IkbIIrQfYocxKhBqB8qVH5BaRmFYRHyHa4r7WQhP2EV53TlYjOhdUQswhCoKY07M6NJpALBrR
OuXAgOgV+yqB2+lFCt42ie8QWNM3JGurdTrAlD+v00gehkTciqVodUot501MfXm1xRH+gbNJvVwW
TnOF1cmo353xZ3F3RRwDhbAPK7c9OXApXpN6aAckunfNOTcRGcgS8SoBrc4+lpnsnhK7q42Bqk6+
fwIU87luXAw7574WS5LbYnEhyUHkGmxqQpFUfqIntIlTNbo0cb5co264nDnw2NAgjKlapJWLRvCV
kqnFWu4ioaXq6XJ0u6rMpBhnhzNVxuXnA3ULslmW/1Bt+IpAJ8CjYOZYesfB0FEboMH7O5yXX9Z9
kZqoKzCSUqLO2voJ9HquKMqfB5DmixtLKq2gecF9q54PedxDhpimSEm18fEL/LtuwFWBGSI22PO5
09n6sPmJOMP/b3DrsY/2OeOvpG07CdswSlwVNfhGmJUGJJdQoOPe0cCsmNfosPnDSHj7YPZqhQjA
F5kBnTg2NQVG4y4AZHZNQ0R1VPcCycEs7fMCImWN63h+Orr7VR72jPZ3y+7nWqIOIAbZXaxS539V
eE3GpBKLoClJNXJZeL4syF8en+0zsqr1bUBSWo2totoWHFs6PnKXtnsijZZCkdesS0rm5v2TSISO
e1FNipFPwM8HwtYjOqkF9YNmzad2FncEkwVL0EzT4xzv+ZKB7tDs9z969Z0tkXNei9u0yk2DaCGd
QLR0Ms7zR2SXi5Q+Oq0RRv9lWLRRUKAkpL5fI61PWQuxRYj7LsLCJpJYGAxmsbeH1u9V1/ehq+TB
69GrQEOUpfMWc+m98tsDsw4Vbcz1iu2DB80eCPT2+tIzMUQ9dLVemoTuu5QeABO5uhDM/qnOKplA
No+82n2V33XKOCPA9ktEUSZ3VJumZbFpK2hCZA1Sa1v/krMjYmL1fOKTQubP+aZ/ZXqumdBQxbKq
vfxFUAy5OYTfqq6nX70JZURAggq77sRq2hin4dTbWPN//hWeZn2PReur8O7vq5pKXqLpC7Yd289I
Ef2Kh+GG0BPxkrrbmVWylQ2OvYhEuDgPd26JIhwtWkB34sxvZCzCfSGM/ngXuE7TEs5T/qSHjS4O
x5+YBVB9lxTVlhU8ddXQw/sNrGYuq06CuronC1E3uEpbg/fqby/VxqSAVyY1Y5n+jwZj515iJmmQ
L67iJxDUpBZS8DBuNkvYYMUcdVS0QHXC92nA8KlRmm6tVOVQvoQ+Zw8SbYoDFQF+8Oagh4yuiaYh
JEMe2g08vijgMZfNz9QWmMabyYS1N8Q7mzuM1gOPlU36aOl7mp9b094S4RKUtpRLHhYJ7kCZengn
Gi96+bH5xqutH/wT+LghmqFEvycuuMemCo3feKWTIhhnfgAtlLtc2Jehyx3kS9RTlWlduKh6iHxq
FUNjvIm9cEo9KecG9UO+kCMExPlVQ1Fk2TJIwoSpcLiq3bq6ulBjuQTB6/MNU5jrpPwAtkE01om1
n1t8gAY5Dj5UXMaGrJN7yczU2pOzx2jW2sPsxBBoP4C48R0GU3gZHghg3ysMgTfaGU9Hf8MHw+oa
ExHtRvnkQ46Xiuy9jPYPTIhEA95piFyMG10fgAcYH6mJel39Fjjg4Ip1ASIDRjt49xNAJcW9IPuO
LYbUMzS0Jc3aTqF9dva52+oBy3q743ci5wzTWxLTcDvBTSTBmwRQhkvNuQNqcHunCg5secSrWDIn
i382iRTTE8eE2t3kpa+b3wJ63F6tgcixisgk/eequuRFbw79MYcdVIHEM3XZkaxikPa/h+e7Zw5B
+UxCsVUSyQB1wKUe9WaxmD8MT46hmxbwMUeF/FMoI07AVlWqhzAuvuZjG/nQNPRDqrJ8dqfDaSvc
L0mPniRB32HvsuedAQ7qO4ekl7GmlamZMMP0vCcxEcxNQmgJbIOrTpXInlgk6wu6anPIDSoAvWgr
2oU/A3SP/JF+zdKiqYHuv3sCtnBYMORkS+tKbdqp/jWqx8qfM++skZxrMHO1dX5ZsfFEZ5huYCau
MCfmgujGd+/QsmBnYMjySrsREVxiXtXRd9YQAsI+nJfmcoslIfqQhodyHgx5cLmfBhgDmDerXfJg
v3g4hVpoYky1e0TtIvlcxp0JFcyT1d9Nmufk/bX3Pf+krKS+lboqavPlrpFA5qT/kiLXqIMFXlOM
wjGCghFC3DC1RBdpxICGoAv+KxryJK87sSHRaoOcDKhb9S3diZHybNjIXCbqsvAIm85JvwKOEXh2
YmC/3jWaPUPJJWf5lhWCyYOZTnPUFrN9O9jm6eUtF24VqzESMlY9Np2Dzdjit3x2htJh56aWOvTo
44VBwhw7kxZeNcMguUEpRerwNG8MbQdSw0H4dX/aITxVaWDe/1jEHahsjj9zoSPDs4CZ7DbWRqfb
jQvV6lg1nu+Xmj/5h/duRMSZMq1i/btxTwFKtCKqxOTrHAiAH0WOMncvQ8pWMJyYpSknkuX5VV44
hRruV0PhTR4JJVAPK0jkvdMI1AMZSceChkKt1Vmb3y7JmfJjpg/9dzsutbk8pVV40+HWGqqhk7MW
IgCNeaqvCQF2OTk39EUjebHyLwSrj8OS3jkYh/ZWifFlkWu4hRRtprB6VkOLNMQ5VNTzd7fn9Unp
ZtNPN1/dvBgfbTQegf+BBz9k3YLFrtrmYQC6foahb9idadqIRP9oxap3yxziDtlvPpnAmeYszXPK
9Ufw+3IuZ9zdPp4o6ktK8NOdWF/TjdsRVemvVPFQvrJLbsOLl5thwXtjZyTLud52xZF51DCfz+Ag
IC3cmaE9ABkgwqNn9NZncG8Obhse/vZ4O+ePt02lj2PnzfhZ8K+G1ZeNRCWHkgIJF733lSdJv13h
nvRhjOvRBDWyRBN7PRY1Dq5fi5XeqNeseXDKcVRwc8zqH0fjdLq178t2cSfQiSW+5CJ4A7Yw+nZf
6WiAc7rSnplPSPfXjzrM6FDiiVegi9sKmVk/2muSjU5wVG+tX9VCKTmPlFYdp56gwCAHQ4z/rGZ1
CtK570RTd4ZiC2ObjynKsNOmjB+DaZkOvZqqbb8Ma1CtewFph2v5c13XKMIZiN+AYO8hs8AgWFC3
yyyZswd0Prtkwzh8o06R2GfaAD+49MDXu93wkq8PBIWz70sPUXmtmNBMZd9MOoQ8N6hiwq8vtick
r1Z59wLpHXZBvNDAqBxAVYm8XmdjTY0JLsgmKcmD/YwLW7xD/+gP5KD31YN6KTDEC0WM+Q1vPnNv
8+6N6NbWon6jxVi5VHfhWvpYY/5ZEZF+Pn/8m3gCa/dYTxvGpqZnfrGxi6uox10r+R+ww/msagg0
Uq+0v+ip624JTUy25AwSbZNZrCicCHwDpMMguEFrVNLGof2xx8YCIZIIfjBFaMC0gZwAb3TVo3/r
AOmCBeYoukVqyG3JUQRlONyyO/hZ3ldn6zNzzXUW9Yqr54vmwyqc0yPl2cSs0uqe0UlBsOXUljb9
RXBbOz48iFNNb7gg1vVQye9sBhggOdPbM/jPUUCt3K389pse7ckkbxmtuptmpk9fQtFMh4g3JStJ
2TEZiY7W1/erpOp3omQd+K2QBZQjZ6xTO582gVTmR2xKQxaHpEEuAqqncFvY1vzKD5aCwIebxZKO
Bn/Y6X6zZ5+b4oyfmtJTAZpoq5zEu1xfbnUfRfPpyXouckZ2Ccaxhv8mA/lJ/tVcyXWdgrXAu7PN
glDJowI3B6+X4DtAXkboA70ct4dcOoqvjGik4WHYj/oc7JE02eq+H+lfvP2GbaR0mjN5bRYL/Ue1
Qs+DDncILEQ1j12ib+1OQsJ2IGFGPV8H9/WqlBe/GOzpbcIYqWfjex3/WruQ1ax6ItwJKxloMo7n
EaEUAuKskSwY/G3bcSm5+PwWRWEMX4IrdBpkMuPbUmaIOWPneXAKDkjl+CT8JiCdmDqpO5KJqJi/
amiznFLtsgRA+m7FBkUr97dsHftouo9k1JRLpxLF24VGzZKR/crdSLjylaZL10/1RI2N4OkxxWs5
dBlT1hUwkjzFqFyg53yL2lj44Rw7kUrrvlKG7Yb+QA/FKo/88v278UH36/jeXqPraz8gBJp88vEg
SWMJnunpe+tR2ET7iTH18YKjcDA7LxWkuNWhtbaYxSnHoZGM0YtIqM+epkLqdS3wG26y+OFWDR2Q
cdJzDTVerD+6Qc8jBBW4JXOtp8WyBCIbEew3Oa+URY/qUN5/Eh7ceftI0OaIEvmlvthEB8TnJ7MF
CcEXwV9t2klOy47kIMgkdfxf3Jiw3A0eVh1ru6fLYiSrIGQBoi3ypat+JnPV0fzeXjz2AlueqhGB
pnyF7kyciKAFVew2WJK6zTB9v644uoWC+Igov/5qMJhH+FnJGdnbRpBMGv22DnY3jpWyULJg5HFb
AUdxyMIumctqQH+a/JjeXOJk0D63DHg58QOd1/ubhT6i3GoRgyUQ+KI6kDezG6Lx3cRn066C5SAZ
nsxcnH53miLXTN4v2Aq4bgQJzRkuusDjPo6oVLjmgd/tL5Ev8D1XWZo6h2OehEppqno+dxbPrj14
j7qARYUWr2MHRjlYrBGjrqeItCD8Wdu6VmcjJ7N+ZCrPFocxozokLOEDsY5qmYgNJiLyRhcLoBGu
blJCI2Rebz9yoAa8Ze+ZFOPwgO+tgSE7gprPVQJUP5hXLdYPAaCAfR01Pno5lFGmqNFnLTaqpGun
ZYE0zMzKYXEAhpLJqDZe+YeokkQGiqK8CACFKkwfD/f504OnmVnbCZffMfB/WtieuWiq2OcHWUCi
jIqW27MCT/f6YpM2bq+1jOaqz8MRhW1gOdO2D+yMcnt3KibTUvRLdziJX/tSvJX36meGyZYgFaEb
5WUGmkdRi+CcsvzzEvIE/GA1r7h+N0W2D6Wdjxqu7z1OwYpfRR5b24s98r6nE1rCc89DlTAiWZ6R
pZLK4QkKM7q+T7KpSBBUfpTYM6D0GZ63ODqJdNWP70GIBs9DJvy/CdlMI2qz8CuorSgJCVxBj7SI
I/7PVJXHQccIlbQmAuxA+fcT8w/DGaWAbjLaYO+nRX+ueviQ6dCZEkYCWhcxChWshPDkCzqDvJld
5wXp+MlwnSAfMWPctnjVvw4riN1bS7S3U6lkjr/upFZtTyW5axVFhubR5SW6k/8uh0FAvMVAobXo
OTeAJ3P2Mukpmk706TySwfl6zX7Den5oL9Dyl5FT3528PU5UTypzvHZp/6LdomwOFIdfQKyqn9ns
wtqYTiu+YKoQGLzRmSo7kOiGP6MBMXqIEgxB1ZYFUHAup180D0d/3KM+03EW2cD3svBZCk9Inpa/
bsyPo3gEK4wQs/Z/SGkUhQUslZrHwqU19k5VnmehS/ErRDsVLjiQtlXmjsKysUYTwZkYtMmm9B6D
6+HLJPxfCLJ2fHQa2GQlYZppXJn50xPzJnNtuG/r/9FZjvXbaoGWjBawVdFTqqbgseVdrqYxN3Ji
+EwEbAPlCLrs10GLO5x9Ovkhxz00+RTG5yhHjkLGgvOw7roqBADTwA0m93oXGmLTJmn+RfTZYrmI
3b9tCxisELeMJ/vgQL2kltSsDasqynFMZYuxitlzw8t9Lrs6Nu3mSIkBIh3W3WYLEugaV1DsIMCY
FnbKyy38DwYdszFeoiX2dC6l/JxJTyBhamyvCv/a//19Ptf5MkASXkD2J+1Q8rl2TfCX0l3lmS7D
Ta6EB5nyQrENWzbBQlaSfIrlfroHY0lAh1GpL9bxQrt/mmxhOUTXbB+SXLwff1Z7coCxbp30i5Ec
y5gOFLuoFZGchKXWkBm0BvTRTOa4oEqkZ7SPsuOIutN8UmKHsDKSmqSH/oMMFwjpKsTYaRngWYor
stsDUQ5i3aJIMzWBBuruX3+3NVD/m5fbtZaSbgS3m3Uv8IqcsEYumtp5kN8pS3+7a4gStdGXpIDo
y5EKi90ys+P8R5bEeKapON19MauBjn3JNaoG7MkCHskAErr+imC4Zr5C7D7hdSg9x05IO/o+pidk
+hiZwE19GS+Tcwy0T2t7xsv8sRIjjYy+EF2IFtpzYgnclqJV94+wOdJ3IHLxUDt1BEAXd9CM60h6
nN5NxwzgyS2vpZ52JhyO8+WBxWKnkAlof6pEZKGaxJJ0QfzoPpjdvrRIwvD5QJGKbTCNMRuQNaVn
extGspJrK9MAyTAYFq9gkUiN8Z4i5Wtjj0QoaYBeWWRpy6fGSXPmjFizijk+b9KHjAi6hPGvjQwG
/znuvWmXHfVjsg1abJ7r57ox8dg3IAux7KuSTFcfJ9podras9Ch5eutFkFE6u3FhDvtEhQRwocC6
sVRXEknltB6cAx7LmIODxYqcX64RxTvRLMG2oQqWCriEU4I4CiGU2wblUygnT3V4tdra2ab5OYAU
sfX+IagMPKjRXj9u62o/4xjXhrs5Uh/AF9JFgAemrDiOrPXVdNsVlb6cSWjwdZYfXyTRCLJ/tjx1
CbDnde1Jmz0aT9VfEreV9fRjwie5OnhHObCGZCXTxbji8EY8mCTKZgn2pNJhzExmCuL7Qw+7CXRI
juEjfOKY1bHVfXEuxz0+ZyXJuKjzhXE6FcJYZxGMo4idTNJ0k2NYEmYpSjX9msm/EYU+H8/6kRF3
2gQPT3s+sXIkOcEp6ihDPnA1sHZkvXqp8t1Mafzygcf7EnmBDj4GmldxtRoFVZq6K9IUgbPZ9Y28
AXWQcEfjt3iPN8MItFqJK6l5qgCs+pDMRPYXYKtT0phjHC8G78IgnK/sUg1oFr/rnXu7UdX/sHOC
uVg7rnSOkliZpSkU76rECQiVu4fNEmCKhBAYqA4IQxsV7hV0ou8FOYqkTpE1VDeUt7tFi++IZX8x
LX3cJEzQYzdB++AaZMXomEYs8sXB+5QwccfVIUL/Pnv7Xs2ddPNeEXFZrprJmrhS8oAwH+JMQDoa
AP0srfLXVciHpXQruU8h4+DPPR2je8798KIf/uslJvEZX6JUiK86BAY8Pm2mhgJJyyfCNyWQPinT
aHQXTs4tRzKQk4JGvsJnvqn98g7bOWiWzRK+FKlu9guZcDnHe0ZnYPnusXAFfZr0d/vlciE/Cx+G
Jd/YsSF9JWZWMRx8WlzesI0mvIDsEIXNF3+mxSlghNWfyGFp+c1d552nWmqcBnP/K9QUg2cIIC+c
12PMi4w3/BfRt4k6hG2qFYgotRi99oWHCp3WekLWyWDXZvttjpRQ7VFnlOj9kUH3gT41lF3YuLAc
U2DoQGcwGiO+CUrLEEuYm3wqM91YIykPLEpWej2lNYT2AmsXpjl22MwgM3SBchQX8m5OdVeRDB+y
TLiqJ3puOuTql07zBmDWGDnRwnh327RSCNw/DVFETw4yrRnz1beF5zNsoLhnxnImhXvx804UW0V9
jEwWC7CbCAAtGKwg719W1c2Pcx0ky2b6wlG8EnpG24Om38HVz7sVzP+TpRQuTHX8E5scogbjiS0l
wwVJ0G8W7suTS6uh1Q4Dgl0wvUrsNLPJaEuD/Cy0dtnw29AtzTSV8PzCNMLhYmQRDWR6JVYn8Azb
TgY2BCoMp4R1QKTfkxBJwxii8Q1alv1g9YRKbX0GWwxkaidcvVue7XZa0fVtXsAp1sgLGSznUBdk
jovM5J3Bunt8idb8S8+efG3cwERx2Skm58JG6SEBiRTr1fuTvrfdcbHrwe/8v/CO16PHaoP/L2M4
oQO3riHWhrdjyF3UzzUR7A+hDfno7h4lrAyGnQQp71uRe04IIzVwSm+xPNDa5WLcglTmK8BcDb/8
0bCy06CdnDpbXetCPHDdo3X8J/9Ap+r/oWb05jZw+Ht/sHgim3etKOSpyXBTFGuL1B4T5COGNzRu
4W+LQy+G+TcuIjmNRvmgesDPAuehZ4BRL/+Xc60GlyV4wQyfTFzrlyP/6WsGp7HYJht9L7FUrVG5
702wqyds6fCmSeH0WwOiIpednrNFPc2zxSB5RiBQH0le3qLCkuHNzrTXxBE6Mp1aPI+CIcPKDUDt
G8qkbm8xiDX6o2KuK9H8DUkJNwZlKKTMQ3hnRsSZ0EKFnZS4RrZfDxunriUM79fo4PudyQ+JUz0K
PGhzFBOXKnPRXriiXxotxnvKQxrngYSszkm9uYVO9DyDn2JAsDMokIVCiqej/rGOOBncv/Gb17SI
I2gY8F5I5DBRnbDDKBxdAPzOsFtBq7hz6lxcxan0UenK07PWI1Olpp7VV1svBX7QXw+5P+reyaLW
93oGgBflIigxEeWQnjOxhjwJ8S0URLT3MyrsxcLdWApRZJ+kCM5HaQmL+2BTIDJUdxQxzYCYNtl0
zBjSLUoCnwZ8J59Biov8SYF74lDuZMZgpRn/t5C8u2NqKzMlXpe3jRrWgWJOHdLAm0QhUsyUaj2U
xF58QtT2KA+uN5BJMkZIQnJ0cG6aM/7//HQPQ/ImV/uaq7Z0735nWu066jnJzZ8nBR2J0F5if1WJ
LYYFR12h+igwihtsDa7na2stX4beDyOuSqrVGUx2EGJQP8ssj8IUbDgeN2lygn//JL8VmKNEnWWa
CqCjBjBXkpdfSEbUBVcuSzRkkle9DtAogUtKWR2GanQmRpAnA4vIiW8AnMRQeFi83kwDvBMAmcEg
6pUel6vldlyz/C0wMcLhODkQYvNuJaylLhzr4/JpsocP9xVPnvXQV/O/zBOLMPxk7g882hUD+VGp
H2vY+7tzdIbNW6F07r7exTisiPS4XyHm7r8/JIGVxra+N76BkN9tChyBBGXI1b7w06O/0KsKQxLd
sT9t1SZhu6i5LQslylVA/GzgbaNXhF6UAKjtCcUymPNx+enyTBfODUUpsqq5RBVTdEEFzHzBW1dm
T/3xhUjqrus+0oIwysapR1UKnIQCdtUN61lEdEACThhirlN0hRWEZrZWBZHcmCgOJxoGLJS1g1iF
a2E6OHOOxCjlS/DnHl34oL8H5QQoDZlI72tqlfsrPFvLFjVw0MDKgvJ1bmH0MrjxEJzzkpPGqIWq
P9jnhqjQZVAXYZFmo+6oatA2YuatwcsnTcnbzXmKXFRJqUrA1KQbMtw2bD+WHqG5ZJbJ34elYLhd
yfKdCiDYtEcP+CGahf7aolY1rAMA1X/+Q2qYMKu5TDazL1GWWNkKo95vEyWt1HyIHsrUcBcUS5Ak
PwVhMPgsrT+npMOPHx1H6wZkZWspmSps2+KnZRutz7b4yUsLZ8yDnDKcInDe3NrtVJ7VHoaq1Cod
P9cHHCY5cvz1g9LnKEb3hL2ZNYAsxa7SNkez7SvElSzsYKW2iASEtSPcfBQeYZ7ZlA7jDJ4Q8BF1
q+WtuQBkzYXIRmDbSkV4GJPrJSpCzG40KPLgEGcXtZIjxxyX9Eqe3BpSqrwnKSwxL65xdEQnlSeS
p/IUXPESnVnCNypudi3ZP/I3jBGPECzxE7RiWhEh5D3vy3mQz8TovOgsdRHIocwQ5kuugcyxcfKP
WHgSnXwDAs1Sc9/RyEk/hPsN2U6z8hsB4cNu+o0WOiMjoVNI7I57ABu+ts5lbUcM7dWPK5NO3jN+
vrl7x6QoZQ4lUIHYpk1jYX9sbiOhGDxHCnnioS8m6oku3OUrGXsAKNhh0OV+9dD7t0Cdb8SZ6cqx
IxHITfdKszT8pHuB5hPnOaly7cb2G2bkm35ht6ySiWbiMOXg9LhlOuhg9Ks+AehHJHt/Qp2D+VvF
UzpNaLsohOaFu2CJDmGdarJv32FhGAlV96iPzs9QczjZl8TbcVJQd5mfYpnhZ0UhNtcnnhhOtQUY
wts9qVN8TG6xcOlq7oHt4tkVouY7dRVCyk3GIi4NlxBip3q8jgVb+sUYjJ1YoD7zUiRzb4n6Vow/
CmQ6IUpEOKlwMynp834jRAWwL8CC+BV/tq4XvVnKfhx8TF+aWyiOSu3kBiwUVW7iWzBHNE7A9yHK
FK+6TwXKfGZxc4eJydK4oYcpT0rqdszKuYqH31tfW+rXFBx1sd8ug0JKCx7b2ZPT+anjmFrYQe1U
OzfTLSegkgOceaTJG1IjOwlu0+rf3AC3WZQDZxGbqGlNOm+pkF+2DU0gJE66LQ0sVb1LZ3VB+vGJ
fjqse7E4i8LBOsH2e0DT9P44bzDglNwaQGr8m/udE5UOJBGiK4GSSe58V8hz/MW/QhVU2ElTe/m2
tAywXbcvAhshEJL89pBMEqYLaFthwkOd8bqSiMzr3EXQuKLaE1GhLi6yDxD58//qxqI8hEfG4Yig
pDAzbVovWjVkDf/eBF7mpizOnXgC4NUFv58TY51xvQV8ldQIKx2kKX1CadeXz3g78ZPzgWCtXAmt
6TxQ5iPS3xU/q93kssF0FPIIBYri/B0VWftxzDibUx5rM6J4me4kCxs8uoBwVaPmcbVN05cB+gIR
3e3mvfjFyXUWZYr4RXUSHldWHeZx94lmR/ocJ8fidKWcRtPT6EYxHZjNGGe31J21mWVlWSMzj43+
qZrfz8UeBKxIxSwBmRMfJX3v6s96GsQNei1jmGybGwZZPNFCzgRGEIv4LkP9Mfod8RFqasy/5clI
eGwHwDwqYHHf33pJl7U0TlzvMm++JQ710a9rNOODzcZOWIqmNNBXXeBw219B7X5Lqp5J1DIFJVPm
wtuhP+J/hdWA0Vf0+rPeamEi7+buJKrkHs7OMsHTeuPC6R/4Zz6cMDNtyWrYGIsms5+10XMw9Xug
CiP2vdpJ92n8jTJ8ZLXzBKBghEcgdDfVCygseSVDQMAQqqHMzvVRGWPlCq11d0wM2hhUbFg5pygI
mgCSPDCUqVBQbh7rhHNY6RgHjg9rZa1GyiD8W4MoBKYByhHbUwGiBLMz2Ija5DPGYWwrvPNk2FmF
TtbNqrBvmkIlvINmCQJFsPNV4vmYYQDXw7lQPaFfeAWGUTMROv3EGCNJ6Nucg4TZuNzDQM93wKW0
9B272m6/ZDvApk3ohwDxYD0tJk5325K5JUqzhp8gTmPeTf057rX8RdDFIXipJO/HdpX+PRX0hcB9
DnuVyoIgGFK+Zh+LvZX8nWQblj66acFCn28xh50xofv+nTOEqJ4AcJtfuMspxUJtBJfE8e8/pb7n
u00PRlnWGmG1IISXEv3uus6o5Gpxg29kNYyIspq/w0tVtt3j31e4RlSisj3mKKQUBpCQiXNNltho
86/r1DkKOVGy7biT06uZUgY3rnTUPP3h7NhPLNZGV2MB/wrrDhN+7on8xYy+Hhtwo9A4z+TuM6S9
z8mIwyUtKB1v5zEhPXjhkytN0rccf55pOFDGJU/tOVmH129+qUCHtqXEHKiQImoAvkRSzf5w9HVi
pmRR8cExhqPSNTx3D7eP+VZiNlQ49aAjy1vumV/IxEi37e7Kvn1WLangOyPoO9V4UJl4q2zDJoro
fWIEJuB7ahYDJKd0+PzoeYFTF5FjDotV/kDhW2A47ZZdycWwikG2GV5/Cgej9pRCADO1NNIf+c1W
pi21EtadWEnR+9/DRJku7Elj+cYltLH1A5MGwGIuQVjPm0TLCIjGRDUj2Dvh+dvpkp4PrfUizMQ+
BtHM3kPy7xaAcpDcJZugjSIY6ojPJYvAYX7VjBdR2Trdv1EU34asuvCMKM2W53NJSj7GE4hXJXAO
IVn7z+Zue7Z/S86gq5CnZsYnvjw3LAZknOYzlzhrso8Alb69aGHt5VfjO0+KIxzcsr0Xfdp81rUz
TTFlLNC5piud2eFeNt+0/nX3+9aCgfYBAM0grGXjnEQ2gJ6T+NLx1LR6meSiR34ozg+8PJIswjdE
i1XkJJuGEO5ChP2RPFM+gSIwQWJj48+3Tp4jzK/kHcC9ue+/B1iQNGYHxMmcUUWUXIeohPXcijl9
NTtAIFlbljcNzRY7xPxpybo3wOyi+zCMF+boRjpMrRaMmDfwgdydriRKZq+agMkdKZlqrfHGQQzc
9PhlBXc/RZU/AiLWBFtCb/1UX711W7FJp/K5D/tETX2AvCHS7nnWycYvoOrwNArJdltmiFz40j/y
YXxnu7Dwx9cDK/zfEcqq1olcGhx1Pk96EP+OYyLNxZLRNAQHiI85rHCkBXZWv80Mmd0uJ/dMzHxj
GrcnVGVQDzJz1sdb2quPw99LF+Syj+3HLo4VxhAY6YkMiUemALigJHHYmDtXJfQ2fqVdL6rsdROK
HS+aSM0S1t3rc9vZG8IlV9kO0qBLo9sAT6/hgl0YYM10BkftlyNhe3044jhYn98X+O4MiApCqKDw
ozzghTFGg76DiLn9K2ZvzQQaTgCPM90PBjvUDvKpLBMx9M5G7zA4o/t1kdJhAdlUZu+PVZRbOdoK
VKG9AOZME71O5/APhLYZg+E25gU3YXVgweXD9XaVxInwT+MnLQUPf4us8soqTCbtqcm7DDT+6g7q
DNkiCS86C0Qn0ax1QJnSbUs6VsbC71mCMDl/9EkjOzyddYnJOSjjTfpsHDnEM89jIwJVzI5Q0ga2
Jr0fNm6iC9SnarAPpLXuXLaH7MhjWcRvF4+bRN/YlgiL8l9i9UseHDOt6AmIsF2HnaKMupBrtYX9
s+a9OdpDManAmBQ3WAEwXohHITiEJVRCLcxRfgoXZg+GXEvIZsxMCUe8fb7l7zbOeH/yjPwsiKHo
ZvsnFpm3c+3YRU4B5OtDoYrwX5mPZakB1gfnbputmGXeE0huIONouNqTUeodXaxdfOD076Y3YgX5
/7yeibFeesM9WRj0Kl+QVuu2G126kteoEZaE+1xNok0slfNA+ZDJeNS8sXDLRAqGay9vazhURi74
BI7p2K279mFgJh5g1NPumSshJzM+LD+/jK4Cgjzuxa1oksJ5DYKG210ONq7nX8aQXjo0Sd0fV2IS
FxJcmTZY++z/CaGp+Sdd/wXdBQWU61OiJV6BwD5FS/qCC+/MKcwUhujPaSwnPDI8UYmxdW+b9sJW
90dTfzKBQEfacrq87RTfvbCNUTmhG2kUm2UzOclBKgPaxWDGYcjv4UCL8JgziZIk26XQXTsvNsmH
TsLNDj34Dt7zcBhPSBL2Hqs4CtV4moDwU2mqX+Yq7Y51l9/XuT1t0dK86jECAykFkpjBh8TAgvs0
R/TNGGCsq/Yn/PwMJErXksreDRPLO+/TM8k9TaCWSc/soEFd95heV1tUx8c/Iu3FLiPPBPlz7Z5w
oqSo4FKTSylFkPffCQ1cl7p5jaBsjXxYeoErw9iP16gHMuDFHQr3fsPkwbhhwHEPdcWtatvZ0px+
RmLGj+uHcPLFaKBcHtfijrTGoxi+GA/PXzH4caHwtPuiSNVLIpEkdFDyCz9p77oHPbZVPlMcva/5
Q2D/ekpjUvrbRV29BeuhLde9yAuY0tZHu5pUYVM3hHqaAsURQe0oTJ3qbQjEWIZGOLQlR9PSCnG8
Vq9rjbIa7LsM2xDHpSWnvxW+Iwsw/GSUgewwiD0bdzWAa4AFOe61qfCrgH5FtJCmt1EXGLHQQA71
g5e/Y45+PpwhQ8wPxgTLt7DJwaicLVJ7j04hEYVFDqSTa+7x2ZNTh9judREa/KzAQwVnqYGlJdfG
HDYuP0dS31lwYNcEW594i75jD1wN6lkvdV3dRZ8kF8RnTHBc4DQ+8ul1yeolkJ7Bld81wEsHCUts
WOraA3JzZohVVR2dgaEvK3LPQQLnSHWYtt8O44N6huYfnzlQaDxS4eK3a/H1MnB7U4FWSq2jTkGx
QxG8/Qnr4yt6KFdFhs36HknBS+3aMg0hCABARPeP3TXWeGbEKP/poCRwppbO3AJcrVZEYdmqVHjv
YswUVEPGCv6t/BaMh0gIgIR5XC28mMT9AO+k0j8KqONLkJUDdeJ7WqzhltofJAX/kbM59YpZYH7L
nsaTpDKHeByS8Xje6SdQSbKkRgpxu5iIl29ayVoUDdLx+JumOS4m94IBPHZPAXMcX+mLEXu9KckI
qXuurZQMqkGsabVta0eCNv460+a0TNHebZ8rromfDk3FaB6DrA+bjKrFWOOKCg1uJzTSVTucBN61
UML3zaV+Ls+w3yX2fUgi7AV2kDjOLd6gRgAtbl+k6QQ0KVS2vINkph+SBiKSkPqOyVgqQSeIC+MY
UJfUPT0e3HysvJwPVXV6Ls+jwjDxO5Z9Hp7fOena64SA2uX5Hbg85kQjMhqPb80vdzL88AMeK7El
PWzWx6HkGLTWgzKeC2kUjz5VkF6DgRKlKKGVdjd37o7IPxBL3tt2HzBD3tBe9xQQlsEwvZUSNadg
z/i49I+NpFGrLwjwVjzwbY2Gkzi/BaEn2DJTUo99K3OI4NwdPNlQkBwgMMBRNXp/fMm1SRxU1hMQ
1VaEX22XL2EOwcK51iP0b5DihpcUFSRaxmlX99WKKuRygffFZUCR1v+0yW3YIjiFuWsJgDflNOj0
VmLb/jof3UdhpuQ8gGxZP0q0tkkECzk8iogkWDHkeW0ky62B1zvSbmz3PebjoHVALai2PwuN3w3v
Yeu9IG1n7j0Hi1bWHdXgTwT5TwH/bWEZsd1H9T1KQqoXGgKSdllJAp0i9V3iPtViZ1Gon2OsmpC5
tlstEvauudRSW5ub7CbVtm9z8gEcyo9nfDt7jjmq7RWHHO5yu1pHBbadEBnOsRJlHbhSsbpfk6sS
pyz4bUSFKGRAob/JeBnDlHFKij8Oy6WFxuxKBZs0gZmou8bjUHJMENH0akaiUbBw3zCEX4TB7zG8
Ub20ithkJj15PHzIjrXvOxJabS2nyfOdwshdrXjbPOfZnUao6E1hE8eqVYbmQ9Ii5+AGWzqFTLC3
u7RmxB9Lq1X8esbcJqOAzKk38UXuajnkKw+lRnFk2+GrObwzPcwL1FnLL4LrdmlGm2UR6tpa7WXM
uiz7MgSxnTaaoHcLi8H/zu9GUPJQ0woYq2itCvZj7o5MTi2PL6C/FNE3KiPyb0klVu1RFFAx+q8a
NKo3iyKRIroQrrX/cmsqI6acY6riGVhMEUzxBk1SUU241cA9a4jDooRYl90uBIibzrInV2xXqDPm
QhdR5wqOoGHNf0q7dNf+gUODFFoMFiOYAO+FlDQP5c7blm5qBg+P1NZ81bHVHKJKd7nRYAZrGZPF
/FA/NDYKDtETvpR3kWW5ddyv3T+4UtnWRMp7EiXavJyELrWyJk74L/VpAsCxl09QBU5viDjY9Usm
rWvJiF3lFyHO998h/3Hwn1o6FfwsyJQGirXI2Ge/D4AZOpUw5q7DD6QD6dJZusUjwmmJbyfJB7lT
hDULLZcXkJ/5bED7+AurlCOVAVvXMGuwbGsSsoxf4hQhx3AnyPJWNBqIMemc+z13Z3hQkbFkrksS
XIDCyODJhx8c4Ym9h0cnZG/L4E+Aby7pD1LLzAjGGkb4e8Id2F8RjtAzYndTXd5pRZOUpgkY0awh
0R1F2IWDZEthaIRDqBg1LjLonFJt5JJtoKOVRbfWyQd7z904YpmaaOVaCilgaPE+9A1+yqTt+Rhp
aaziEwP7AHXAEK4ilzNlSPtNAWAcSQyHBp3DpkeT9gvQI9W6lcn9d4oOMcletRgrcoAlAtJmG77s
vLQKXnXzlyPF7YqiZusMvzU2R98cvr68EiWXuAVw4vm8hBUu5I6J1TIZeQ8KnuZtrStX4Yc9d7h5
gLM0z/ER0IIH5tqmCfTrIRkoD8D/LhZkRlLSqNdwlXMvas4qGJHTJ/pP2aFgzl5eRWGqM6tPuXFW
L6y+bTdd/XrYQ8W++wkCPlBfVlaCD16gPymbCUt3gc1aCzHOc4Vr13wqPLlMC1IFkCw4kWmdVYf5
EJIhGp5pe5GoeL5KgYJvaxTM6W5MRZY3Hs3xPYg+od+8NaDrF3tt5PnOIPUTCRKT1UXJM3zenDg/
a9ZGcnbM7PZwsiNt2pNhD+lEqpM3im6Czf5tbRPXjQJyRNrvAMTNYjokSS7Z6Q3YuuMz9vM/KWdh
emluJj6yJTc3U59Br1FNCa0MzI7R/knSRNPyTNLAWIy9O6dr7xhEpgdgeM/Cgd8nnwB6Mg+yeW4/
b/s8i9l8MuIUx/NL3MGKalpzMSdqc3awuw0f3+Szhrp9DqbaRowYaa6VQeuaE4wLYzQ+7uh1ACNd
8YUcdAPdDzLmGdolUoTp6STlQAnAaTpZ2eUz69ITHWd0m4MWRUkOKxdImQqLriUe70ZD4fKAxw6b
dIB2uMaQ9LRqYmn2FSQsdiIPGwG5BjCTdMw8pzvO3M6MJheKQb7JwWtvCGir10RRnEWdiw5xiDEn
OZl4onx/uPToPjPsjwyMbNZJHZSj3BymdlWdzzj35qrg4mBuGgBCFtswMDY4bxfH0JndVpEbT0so
BPCJ+dD4bneygLwnX3P3p3VYCjO0UPKQUGpMcSRGc/I9L4kuk8rCYETfAuhbvq++/JMLr91k4I4l
ehofhnLD50EulXyvPIf5EdjnyYz79K+n7Cyct7W8P3aGQ8GokuCBlv/aNQk0hBXPxbKg9xWPyxC5
wlGnkeHp1FEVI/C7Le/qoSy/tsuJ6awfpRm5ViB2X2sLJeyBJ1uGBmBgpzCyNvHurlqMBG0Q5Clb
k13xuIcOHpDJMquq+uXiXo0/ngTu+Ug6wpCBeYBL0TuSRDMkVOjzJZiBQ3C6DQSbEt/l8tQwsnAg
N3fiz1dhVlJ+9/yoaY7m656e5h/kN1Zv+F9+71v1OjT0ZZfeEYw9NnQappqDRKxuN7zyX4kQv8V1
YRS+YVNY9DVyuFjYkt19TGv5jmMvHXWtgXAzIm3jpiqWTBvGSwJzJuYLiXv1u19yJBuy3HSjT7tz
b5v0xHtKRMd0NrMF9JgDKTkIJw0NThnKfqsq2fS8go+hWT5ECV392tFRwvA7hvJsPuBYH3irJ5Pc
vFeyQeWrx3f9k3SgOOtl6C78HaCBt5eXCowFejQAm4nZWI3LewEMc75NlhcXfNGhDTPzx8AJ7GsX
7l5L/UGjuhpqqJoJWvQKeNeX66ef9pAd1XBVn/RhKOjvK3DlZl8uhU0MlyF4LkMptHZx1jiKzQ6+
vPs+zpEcnNLFIDGjJJpXKydrZnGIz1Je3c54COrmZf+3wWJFF4PesWH9RterCRzCJrnH7gNBMlti
m9Xlb3drPwW9242Rdx8ScwdxDMc71yC04kjkhLPck7f5W1+gSwLy/cdGkpz2EeQW/2jj6edHuoVE
PN/litPI/5PMvT3olLPeKW7EAd2dUSTvT3QxrvyDfMUfJU9NVm3wRwWIG00uo5Dk02cpK4SGpgTo
LkecCQ4f2k0g7IInH0GT3OjtR7KKUaCOjpe+R34dAuiq45arIeu9EP98zvKW88c/UhKiVtiycKRm
/nfgUzRAf/0Dhhg00aohqda7+4ubOvZsusBqzLk60YNiThAvb1GgyBVl4iGdhSropXcH9oEpYPam
6oENPIXtHWRN/Mh0zyxGMThQBM+urqqhu/CGGfw1gx4rGVmSe/LkVzxRQ7o3Nn58zEyMcbvPTB6K
sXyg9giTgPLSWkvh887dS2noLiRNKtsc7GXAc+EZmpzfuqt/JXldwFCbVchldtw38JicVUq1TfB/
MqJvnI/4Parhu7sKPlHJYLBLzLxpYnAUnMiJOCnnhJzn1alTmCC+PmFqNDQsdRtzoUUJayBzcmwX
qNfG4k5V0IZeM4GMvOn+sCaWxgcUmnXp/gwrN20KnkhFNisLXgzg31dEVfIb+KoocnkSjZ0CSy6c
kjqRQV+y1NkFB30aN5eDKqmlFdOP9rt5F7oSClts6sAArJF8M58WEB+e6mq/QvGshgXeY3sOVyV5
8BVERYeVHKZ32fNze+tUoA7rdHZCCZSQcP9CweepBUAhC46gobhHIzCeR0BdKKlQcVtxjO3cYWJr
I5VpR4UHnkktyRv69QNGy0hGqwZz+8D/vteFkRciH9pa9eP/CBjC3FVou/tLxzhZCLaSRTfB/fi1
Qmut2EJbh/pgMMEEnSH00vVEbywPbjifE65QP29p4PfAEIoeXAjuAV2vX9v0ol4HC4URIoF7vza1
yNRqRcxpffWcNMGIq1+oZqCKPxWD+oA1Hng+ZJN20MtFL0P2YfaHM3OOrT3jqtBRbVJfwZFhCkBQ
nvU2PVOIUDQApE8JOGrMV4JeahXdwWqIhJiE3M1blerkzsu9oV8+83Y6uW0MNEbZ2BKVwCmGH/6p
1fajfn1sYOuFZr10uRCjRDlr7M4cnA0nKO6Gvgz6O5iPIP3qEbe6Kze8gR5OoQ6PlPCdR0m0TRsY
XfaiAD+geJ0tXpTMoYhDCW25Gp9pLcn8jeOjBO2HMCBQ+5K8S1nCui5o0EPmi1X51qiZO862/xUc
7ao1jFf/cGYSDZ2BDmwDIXDt7ZVSFbVyZYG37lSUeskUY7PLirUMKppAbX3ZfSKbo0mXorA/+w9N
LCPdkYy8tk5urQ2zzAvRupZnGXt/kRSCQjBffk8KXo6riNExCH0VeSxLSmCLHg43CyhLusWaG01T
kmOTUq0/iv4q7PEqcUq9ethqT06MIdhkhh9u5WGAV5FVvH/3cv1sspb0nxGgZrU5V50yUCcWPa3w
GPuPpoG6B5pTVD/a3PKQbTuNt6VTVGE63qnqvkRDUBlM9rYb9rU8SOINiWD3hn3M+CbFXGYJ1VWy
yIhzcmXKXbCU3S32uK9YZR1HvouNwbiysk4sV0zCaAxGwcJQXpoqV60AQqcOQ2xDvBeGN8sf4NPl
s6Z9FQY1CFlKfKeZfQ4Gsr93dQkOVs2DrH/5ktTivGu6yxILUw4U0/3kM5QrQo38hIKqbKQ302ON
1sV+StwDMmnTc0hI6YWYX/CQpvVVkrFOLUURewdfJ5Qzp8PeWOJty/zreDENrUzsUoFdS4fC+Gp6
3L41xnarE9Accp525nXekaTJzGtbPizuo5s58jNj93LrY5MxxLTyDLsd23oUAn7gVQybk3bRd3Gy
H7ENIacw3g8TJHxX+NGLnnx9rE2oUXQIY6Hhwvvpucx9qCXqClEGZmk+Ai/W/IPw4lp5UPF6q/Xj
5nmt2r/OPZO3I9YsR5Oj2+/r8IPxUceQ/KBohlxcVMzDEf0MSpRkOOp0N/b64gVHRcxgP+F7wzPr
BclSSzt9XGGd9JNAMRmWtgMFiKsEeiEnaMa2QAUiFUgdZ9mvF1nRQbCZvHHctt9r1grHxybaJG+F
0WCmh+PwYHdo9ULHL1Riz6M0svfOlJd7zaHDAamTvW4bhHpDipskfa64CMcSsP3sY3sXMFsxRd6N
7lZ20gkTDCIp/VObTEjPFAjXj1zmDB178DHmGk0icDnu633wM/4r/630ElQCCkJEJ1f//1p49aSU
D1yPMI+GzKLY1M4TLVHaTy06AF9ez17M+dHbm5JLI/hz5MDX4F87DJk7XZhZ0ITbajSumqf88ez/
IJo2VkS3ETJr6Xp6UU5tw8UZ1/KLQtrUjiEUaVTRFqlMUt+NZmKOQdcQoXfd8rnX7uic24mUoxFb
xP1FvzqU7qy67CXt0ONdzlxFonDc0yx+gyObqueRelWIr9hdYuDMdsIQ9Qf7WvhpIsO8nmsR4BMQ
ST/GBxlrf842THS+t9LNL6N+CFbUVChfWQJ4xvVFW8pEf2KhnbaYaRoKY7rDVIOp2+P3COGmSl6L
NxqHtTrpdIu3bRYl6Ph6ZuAKlro5W99BZQutkGJx3CvJOVw41P4eqjEjgWxnfl/P4mOeXwwksjAz
lPUrmE81WRAKoUzZU4cuSUGoOt/6qtUlmubkknpmAOs+nwp+D7E8uxKAYI256U4RIAsAfYRJuw5c
J4LYKL4y7iihQgg6HMFG7NrWcbfggxx/khPDgBqdoxfZMsycUxIPXx+omRkm8GWvC6LW9KwcllXq
XCSztURkyVZpWFiA2cO4qiu9sPDn7g8ijVUpx0l6lrUHYiNZfnKidDVtmciEgurPT6auwsr/WXqb
UUYtR5Kf/f2gzx0PHY7Yhhkrxfz3vMw3VhbkPiNQOQqkMS60FZaDhG3iCjgokMUzS/A+EYwpDuxa
vXIXO/tdMGsV4tPyBUZcy5ufBWfUWlYbeC2Q5zWICvwh6EO+vK0kZ1qcILYMLIjNQbY8tPDvP6xb
AUc1OzpTP1bXEOWS9yE+OVU/Q2GKpYJo4WHT0ItDjPEeN87RUHUg8wWsypH4Hj/guq6dXFBM3oVt
JPjSx3jvPRCmT6HT0OlDV0RZHc6iK6BtsVLsoKpKMKaV9w/tmqf5/kPwEnKN+9ipUSTj11s1u+jM
gul/NcSfUO4m48Zc5nEUbi3dFLk/r5KIAsia6rCjR6wLwrAXw9m5Cw8553+fGjlpWliSpBmwCv41
sJc2poU3cIUQ8iUjmBSixKkcppaYsQnhHS1cnG1af1HlRpLjSfkvSYpxuMakJj2SLVXTsS8Kk2n5
m4Y9vt3kV3YK7etyA+PiSwlq+iT2+j7N/PaB8mfUifCZQfb+xV+eZd/xbNR4WYqsqZB2RPH3VdIU
FyGR1lbTDceuHmthf9WvB5e/uPlV7/NNKH0m5NGLEqr15zkak9Ans1Hy2hG7Hu0WohahjJZiajPH
OQnlIp0rlaYdH/S9ruhIyeodHh+79LzRiy5si5pjSNEuyhC6Ch1SFOwnB4IDhDtfMoiZ0hQHVS2M
OMNd9PsUz3dnV87Ea608VdE3kHeO9FHZvXJc17x9h2xSjUnQqkOLiSlZD4YCom02QHuKM97yRp8Q
4SpD1r6gP8piaiRVV8OwkMkR06NBx9ls0lcuH5MPDkSBCdqLwOez08W6LpGid4X0sADsuowKLaLe
NPy3pZfx+bx+iilJPQEu6BHylVSHmTxcxg4/m9Zs0/mzgTvp0gNBYjI84KmnxD+tWMqsEtgU89Yz
SsLJZ3sWKLfoWBLzdhNadxIaDyZgirytwrHI86KlzNhTK97dnPNHhgT+vvIKzLW2BrPenRbsA3V3
Nr/vOXG46+GSH1VE/JHEjhmrlw4T080wQag2AfTlfb3UEN58m4Dfeyq8ftohk1APEJ8ELnUp4G9f
SHGuVTxgWVTSmbsENktZL6xux3WMmY4U0rQ/vgIk1UCihEDC1lWQZ1sk1FXqE07dejlCHq9qLjYh
tad+Syw55dMFrsUaVqQBKu0KpP0LP22xd6QbB8iikFreY95RD1ui4EpFMmqk/YCs1s94ac+XwJ3/
a0xh7VsDoo2pm9MVhymAAWcbX0HHVs30g9wvjzOT9fLr5E2XToecX7MzNKOiPutJZiixrjEOgbjC
6a+py9sm6ygl14SP1pETd1a53FKrFOZtZtBt4pk02vSKgXyHMc/131w+khhPfRO14hjG0apULcEI
BbmX+IWtHSZoSPHqeoBhLgWf3k0dtqZXGCB7mf4sgt48qd8QupVlTy+OF2ZMjKABSyB/fQO+fLE3
a/g8IMwId55+vmmia7ttKioLBq0clHh8wZWGZgbtl0a+/T9H4SD0/kiEERAo58YW5XDjr7KlIEht
XXbZrXxpQiEanZ8RQTDZmRmVQXXekmdDDDkKqV+vN5eFiRJEDvtn5M1qukcca6sBABWf3Tt4CNYV
eyIualaGa3Yj1lXquMVINpCPtP2lXwRII/b5Sy9ciMT//BcrMuauKf2E69JjHk5+JamYWbaON3gn
lXGKtmMnCcctOeiC6MnQwr3/DJAXXmaLVVY8aIjhaMmh7VEJUhPkMrUbgZSm45MMC49EePVO0SwY
06DboojpvPOJ5OtP1gYOAnSbH8x6OrZs9PY=
`pragma protect end_protected
