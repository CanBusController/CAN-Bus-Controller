// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
YiqfbY5YpYimf3ryEFt2SlH+9NzMhZi/q3OK2iqZ4sSIaptO14f4e2vE4p4COCzmFtkUdcRZ9SVM
mvgNLMneJm04P77gvBpm/ojuhY9fclFtLZjCAEY6aSOqlvtrRBHAtCNa3W+3yS9Fqe0JUJzfn+7f
TJMRWT1Dt44VdXkFJTkQm88WX7e7uxNOV4h5sGfnVk9CLkiwq2Zk9cDO9rSg0n5abrULlW5c++E6
a+idR/rHCLsU6sO5zIPNZfEIRoYwF38TdgkjxTmP1OmtGq6mDVylpPUP34x4N15zR6PVWTW9T4Pp
QkxNo5yupTVBjSHNNaXj+wWuLoDI5/xgaE5IHA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
O7HFJjr70B12ma/pX5W+JGqqdUpz/KRfcG6BNhW4tANBfDACtjkuh6zUthJEZ7Y/kZ5GiriB2eEV
HSA6I53ok2RoxtYX3IsnKSc34S1G6ZbJDRrl1n4XNvso39n2Cma8dk/0AkbMUxmhz+D5crfeKxCH
ZH/CKmgFmpq5xEYtGYlndEXi67FVp+6C3IHfU2SbGFF9wAz+4344QeWYwqDurySh0UsVIe0g36Ch
gk2l1ZSBcJRkWgm6S4R43MFCeEdDj0pQiDKE8xfTBQzCJSYnA8pfUe86OXhBRybNBHbZwz+8J0Hk
j5wlh/31k+Fn10WQDq2Q9LUuREKuOdGtgCahifrN2jmRHm+Msw/S5kmiAYGxJjGXvdWgVYijR2Pq
yBQl1snBCpTFMHYyaf90gnEvtsgBQHYTE52LuaFSJmGZljIVlt7tNjnkWUUGCSqFWco+dVcfb7GE
rYA3xQLxTTHAGN9q1U82WesB9/fa8CFqy5Agj30XIHerZwEAntUFwYg2ocGLz6jKuC55BxqIYny7
rYgcol9UbI8WY+aeIyNygABvA+/lrN3NmmsUeywBd6JmMVHXBQ1EP1uGq3HwajWVJzrTiaJYG5j9
Ma5XGc95VAqU4oATurMDDdZgigUkcjxnF/kBKkAR+HLUXHpXIZvd3Pj1rDlreF06OYCU1OVxbOvB
4qpPXY4j1Wte9g0FyuYolYThJcs1I58rY06qRH97n5fwSuPB7aInpxvhC/w6reRWlmxGELNKPCzB
6P07j4dlPHl8pZd/JTdW4gsltoWTyWfFboRZQ/6BX38cqVLVdP61sa5eKunRbOBsx0vyvbhSHiWa
y1POsYV4aOrUgPW7i6jqyRQyrFZodLrQFRISk5tKPJb4EtCuHQWg1IrYME3/PQycJe2v2ODWbHld
cxmtrQbX+GT8VKvUZgSBbKjNEeyADjRJpiiTVHgQg5N3jdJqKYuEz4L3Wo41Xkrh37exSrhjwuAi
gz6rQwY9/jdVzsIfiQR07k0RUFBGEdHb5W2RNdC3t/06bAaRA1DLbZMiAUv0hL19r9tUCRurMvY/
uvJlBp7oap+s8/86H+v1fhhe+U5jATkcJOmZovWYDUwpR8Ovx9JLswNtaUGlVy4658Qi6rssbaL8
Dcl2takn/2derKtSsrjBHzKUdPP25Dya/pdAa/JNgxTEhmzDF+2I4j8mLKybsmi8JfYQG5X0Q9hy
RWFKipuzq5aEpFAUzOexPjq8lbOgpxlhjawYg3RdvhAalyLJpaPH2PdhuHKehN8OqxxMfFnWg3kJ
wCfdwv1h/u7lwETAE2WuqG6CZhDQ260lXZI7nMoZrtU/JsFsmoqMFvUNlDUFUou/R0HYn43bqdqa
DYybdtO7KjwNsUk1m0EfuTbtQAkHFJKerv/vNK/IqoXC4/LSt+IvExNKPUyzhl37l5WfyLEgOn2G
SqIbZKT3BMXwQwyi3dGpRmbNI0sTum8eiPaiGOEOzkoAjTfNTac9e/9/5ZDYwT7EaSNuCpKT81R6
07gqUAQ0pjdsPJkoI87Nc+q4O7btXw5ijQkCb9ecBda9+ecG1KvAB0uqB8ccS9N2pNlUv+b+wBcv
hB6onLYbZLQu8Oo493ocH9IPXXnroEaPQpO4HGo+gvpshVwX7MVrH5VWgGKMqdlz1GYtU932SDMf
FHfgyBgFB+iedBjT9KENmCe3lxqnukZ7r3foKeJQ9p1Dyl4sS8JB0EFrcGEaZLrrj6yYDRZmbXah
GfyVstTCHWXGjJ8Sn+Gdf2Y+625JxM8AlqVCH4ILTz8HNFfF1jr31mDVSpE6NXmNnQJ18Z8sMu2g
Aydy5mL6S6LFMcKyL6wRREQiHP+Y4N5tOm9U4EUqkbJ4BIm27VZcJm42lbZa1do8Gixk/QiLwltt
tWtd6BvzVDy3BEwxu8PtD7TYWrmekywfyKZT7D+sai/0Uitu7K8C0vJ0oQQp4DIYB7+FWtE6jScV
1qw7/ajBeQtDYVgAfUjnl1dsMPPJGr5E2jmYsdaTmJ2BhAZiDwRuZQcUPQBJJemHDKhIuZ4dX3J2
FWN7ZawXmA8TRjm9UdkVGvUVUgo8x7A2f6/Rsfc6d3fGOh2zlF9r2hvj6wmSPkZC0uXkLfEJbGli
tL3INvxJOt+l3/qhnZjAV2B2n2++gGsorT/lWj+tkPaEWmW3+MZsWM+1MedxIDaB3kWytG7/yP0Y
2xlWpW02LJoaxHaeOALnCES+AvhtVcy/N33X2juc6mJxUNiWKVIoZImPINVrC9g9a05gCvbIJgTW
NSNuiI18fXWcORpo/zjX6V91T7kMMCbeYc77SZq2I1d7AdJtU+2OlIUF5SY/xsYOgsKtB8wbbhU4
5DkEdXMUv5AoJLaRQIzHl7G3F2aigk7Cwk+PBPU/SDEJnoUlM20YwEBnsKtnFKIy2V6XACqX1mwq
jEr4CC7lbO4rX7EO8SO+8LmM2AE1Z07315dZ8Hg5w0BfCN8m2bw/KkDGzIHEt6Tt/Jthz1Ovz+gH
Na0foPMUh+GNnSfmquWZBFP31UEkw5BBNGtO3TlXUuRaPAkgtnOJBrGtofibCxsQHlMVY4Aihcgg
BIGAkt27jWnnFdkYI7Is6BwAuYNLt2ItOLnl9dK+BI2JCSPel1wbsKhJLtJ/UW7p1ZBddR+4LGr7
hoHxWjOL9OyysHYtkHTL001pHf7tHkcVBdI/7So5atNaNlNHaKuwYefTY61Hbk3ewohx9AHEVABS
eAZEdN2s5KRcS5F3ZihsKSck182D5EeFC319xMQEOxZ/8gR6Se1UBK8Hbh6jpzlfHSJ+LAsewkVC
v8C+7/8/Zxozm06KpJKVsub8RDHHrIlrKgAqk0Tb/XL++dbvi3i5eom4KORbOKSgSbbjrk9eZb3I
1hAC1ZSxt/RAutMfjcck438UrZkSc5/5SyU6PXcuDxJCKUKOQbFbsniqMUm39MRmDafW2H5HCTiN
FMcoZNl7EdM02FL1uo8C1VifwBHxFH2dfj8ZbT0A6KNH92e411KA9pn2WTMiduQOi0Q/yux4+ncI
nFFUW949msdHTGFFdLSOzkJw2YV9R6eM6lstpBWBtG2gmhsimIz+FgDarO5PwfKolbYyEm7tlnFJ
hnYcRGQvy0LMOoZwKF3VtUuNLq+IX/qSG91blYE/lOw2/uxG0s08n3vodmj1vrmyB0MAGE0H0HbF
xTwwbCdkge+mV97Y8r//xCrHmu1xuis9rnTbp82t95JMoYTstlfZoEsmskPsWm5yxrH362rUrLR8
taD+61QtAq1ydszAHLXcAUEPXkoX7/ZB/4ieMHPmM2LhLdcidYd3zB9FzsZEDx51bOSEiPvV77wb
jv5slhbKbhdCal5w3SZjH/hNpK5kATOAgLt0VoMfSqusczI/heLbzWOCel+t6qe2AnuKB505AAuG
liRWIrRgRhfvVleE/Alc15mBZhyaVRXPSNuM8oIPtLKl1QXIzB91+1EjZ6//NQWy+RFcC7TYH03N
TiW+Unq7/JrrKAKN1nynSUM5sZsDwukc8p2LsGYka92s4WsBvE/160hIJh7iktldg+4SDthwr7d6
H6CJwxVsfXRd8/7uviPRAVvu/R0OTWSHgNhAA80oN6rgq1T2mNaYlr4CBCSy5QtvbX1TGW5OK9G5
vHAxnE1hMS97qhpUL5l/Gewo+LoiTsIbUdkRhbNLkDsP6M/83z4UZe19ijDsoLFqeJornwfRW0Lj
CGkYCxr0oocSGePQ80FjrvaJrzFIlFFjoU9rlv60xbAKj1/pnVLjhgmwSmgjAIk1k3Ne4R11edby
rdk1+shtl4nu1Q3nOID6jptvO+EX5naxZYV9DzMF+mG3bPZzaPJKLZNscm1+uI27h73rl8/zTYrx
pSwzWsCr3BkSF8wnSUchWhBaLTUR6q08WwpDm8Rn3IxUnqw5elUph2TWq92r22GKITcFOVRDOxXG
XfQUj6hkg5kzD2XhLxGhQRKiA1Ky7xWfBCxSsjfyW/tytOG569GH1JrCrX+K+sFdjja/5WDv3d48
8l3cPZFLec3xCEzWVmxHL47wd9VP5cZ8nFoG2hKVO+wtk2Fysjg5gsWmonrPFwtmW+zQZvktRBc/
hT8K5dhkQ2sYYvETX8hnwAKxIb2BbPgNlN9oQ9Uz5fGYdEDef4uQeafrrY2tgsX7b82y3v4edT80
G3EQLB6G/e8iTKzNHFv4BbZOOFzewH38Ph2MXMeCHInSjY+t6SNrCY7DhaJn2nfvUqOGx6fCcv09
hj4y1v7M09pSmtCYqTAcLHpbxderFwuDgblHO8uQOtikUgFHLE9h2mcQEMGKfuO3j5vqXkZ5PWek
brAz3weVaLn/IgqTVVzgaUgIohRyQ1E6z7m2q21Zdmp0dl7qI6Sin2FMxETzbYbf3L+LcppJjTgU
jGbepcXdzp/uQemSUIsThWQ29gEwZZwTHPbcvzYLjK92FS8yLtFw0xjr1xB1s5cna4dmLr1O5yuK
72lg+Opkgjq0aAGednHmV0i1PSG5evfFoLiy9e/8idcLYL0bYygLW5ZQ6XaTrXs/ttJLlLKIB6Ap
ZjWtea7HJMZ3od2j+zqHdVCW7ewbVroKWnG0uG4SOoNZmHUHx0lXyjfixc3o6HS7oquoM2H3L+nC
XdSSp2itmPPtmea3piflrvjVqrkaOTYq+hyOdzpKUCD61j9xiOrEU/4X+WjZ5udJQ/be5K3ouML3
z+LYuLZlrZux4NwWrWgkDYKFap2BZhTE7VyAlG9z5y0mwfCi4rj9ypRkKwufRwn9ZOLVmXcfBbAG
HzadNS3y1EoA5dPJ9BgrzyI0YTF8JucdY9HkqP45/Gvzo4hoHGJtYXXfTtwrcrfI+GFDg6EyYvYA
CpMr3P5DQ53iOw/VorD+sT2EzM1aG9SzYApva+//eGiY1Vxyi18AmprUrGjauYXoJkxhOKLoJgI1
7OEwj/W4lA9diVdOPMd3VBwiWSQRSBRQQApeBT2h/9tEO3jnHtgWyjDO3Q/D+W622DIcEKBhfyak
VsWD3dL4XSvrwJ7bMFE6t6nniN1zzSfIHnbzdefpD1gPamrYCoGzBh4/ZRJoBudmnYmowgG4PaSH
Gz4gZ9n+Ghj3W7mwbd5Lb1u4HBfG2IXpbnFtsBVTEyedKdhhvaoYNWgYMF9L++CgZjI5D/aiN7qM
9Mkv2BaxbTTCrX9virfftNCa9abBNum7Fvvs3twFBEiiWqFXX1IiQ+6axsnhQaFRs+lbqXzNxm3Q
7sk7n5H+ZTq2jYncH9vtJ8dSJMMvmXbaHSrBsH7pxkS9OB5aO/PLF+FjNpCW/czaEPqu9/zvHOvM
jMKb9QUvZGZGlT1MCffAV3NAEC9p4I7X4V7QQPPtK5P+KwSjYAE9uMTVVh5Ni1Tj7nWJqKDdypmY
VYNEVkEtgkIS3fMhScVBKz8ecOb5YyDXgwBEkPEam68PSH+Umn/fXItk50jqasOCnJu8MeId66t4
ybuy7fzm6Ci7S9dGgiwsu/Wa51zDFnQwFDLSqKzt8wG2OVKXuOtXHwYD9DLf9WOntuUbz4ZuM5Db
cRchJ00DSIiOoMQm+/wwMiCcS6sTVadgWEglfVFAykdmM5vqG0bET9WSmtnOOWxVDlZUFyYLjz3M
s8LF86l9kehqIPK67Op3r5lHr44nqYecfIDwlf8U/DRHoAmXD/ijeoGGly3dERPqg/p57sY7c4he
YTx9bld09qJkqB3APbeY9sv9UWic5uqJv5N/Vm2roBcfesm2n39bBNjL5x18kUCMtwP6ivRonro8
q8mEuHVgZVy20Tv3Fx2VEmWVzg0hebakRHV7KSmL2OF38g0JXOkiU+NZxiUjOH5urSnXLzSCIcZK
c4Q6um9xU4aixDzmBQWjChyoCgGQU8KOaKHW8a42QXKHkbgvEzBXMB1aEYKcCNGs23loGPJr5Eik
rfi7J+IUBXYM56Xq5Gu5kpL8ouo3Pjo4d3x/D5RTj7CQ01c8lQL0aM/iVsw8P52ZYHEpDNH+6dXm
aoJn1SFg8qnb7N7/AF0oeO5La/aRaE+ZrWBTYIOt9qYC7Ru1cU3PrWViLrQz7B/tNoj2SnYzRWm+
Tjio+EZRp9HPozI5XowvM/O8FE4nS8WWj/hNekvG9QMCiYIVWkj+wGDfJbXxQ64bndWYy/xDj2oh
Q3iTRpDcEi3vCu+3tLKVEEuiS2R474lxTDtSZlJ91mMCm4aGC1lk2rRyjEOscOFfYpI+3oN3jyup
5B2ZWcQRUkpxZR9gmhfhRzrrCUXDsMBPfvhmBx3Cfl0QTCGY7Hi2HaY7EaNEorKVBxM6ir1M100Z
ThH6y4d/nkpp1hqZtKpaxy36czcYMdes7W18CyMid8lNwxCUhkcKNCmoolBLKUX9jfAzxVaW4oRY
PU+bFsKZ+nChweoAWj3pG+8/i3DqTxZBNHxaE3eFmFx1mw/mhKB6SAar7Zj7ENtSNOP1QKUUkkB0
yc0godC7rejfmU/URLKCoO+/GTJMXEzsTQ4T1C+j6jEubXrsVH7tdrGJ5NHcyNyxQvxNJOoRecSQ
N4Y1qGrT87AxjRasce9ttjkt3nn0e/FYaVTQ0W5qD0YhPk25BYoKmjZlONjSHhhVrWZLDCOJoEjC
3t4ymw0ov9gUca6xyoZYbi95tHWGXyf8loCj9UGtOxqcbD4SP26R805e8X9+alCozNSdQ9IFzoYh
QhmYVcVenEoY6zXg6Mckcw7pkSVcUB+0Z3mu01PwhQBwSU26N9yeqOE1gKalG+FLucZW5bd6sZyn
GoMkWXo8/MASiMkZaZO+18ATkP8dAFbBHgAKg9TWZSzu9sRZYF8rxmSsKtVB4XECCIEifL40Spgq
4oiBQp0IUiXJmHgU8saGupnaLqx4B42GZyt9t9t1xIai6fsIrYOp/MPkLn24Xo6Ash93CztX4UmR
0iZ3atWwcHMx7OCSPc1J+tEnfOELmdoS0mmrsMOjju+kpLqSdjyuHv0liyyjmzDtGfr6Yg7QBfoq
wbltHMUT8K5KX389rbhvJhPn+1qhp1bhTPBqDWkvaTRa8DrWUiX4ovKndknzzQlGB+dRGrYa0o3Q
xs1moo7rEfUWS8jBx1hm8bIN0UZ9tz+3OD1gwdqN7FCTqW6Wtdk+17PsPLM1xJo3SOVzELrZDqLc
9vn8JFqsURWuQrZclUDdrOWct1Zt8CfC7RNQ905So4XoO1f049rJj7RSyM9bQPfowWZCtEzae6+Q
BVcSEcd04QRDNQCcufMzbBiTr7jvKwgI2w3mBCFPOIWyM9UYh+HGCrODicW6UPHKxq5KOE2uCSet
5qjudMqoM4TIhNeSc2ELTdcK55GdbmiCBs+8dLLiGDkwA9DJ8e/NZvtrcyreNQsV1DeaK8bgDn/c
lFxWaknzhri8FFX+IHbmr3kPi2FPx3XuwcU9NpWnVOGS/BnqE6h1f3/Zt9pGFgY07sG9NUHlkhJl
vt4hH8qSJwlTIy6uGWRfbAYmPYBK61OyNEyKn7lrhdZNvepWEWOIlaIrsizsEFW6zpkbzwdzG6y1
eCJBWvwpe2QhhfQY8KbHH6EidbrmmGapV71088sNIbie/aEc5kV2HbdPWGJlCUGCBfhHztZN2OjK
Jjq1A8SKYlMa6aRrCWxcn+IDya+AAK4yT0RwVGyKFH9MAkntXTSXVC9AqhCvwCkePYTLKpy8/74u
Xhi9VlxAoKEaMgawf4Znhei/QKDiBKi46I4Nch7ma5uQ0bPIBKGwkSNq8Tru8+GU+iSBYWSLcuJI
wCmegIMEzri3GkaprCOpdhfMFFgQdqp8Bn7ewmtrsKEiO5u8i5dPayWEgm0SdKwJFwVHslXOEvbe
4YMPpok098dAoeBHg0w5ExLydmtt9bAhAz1JCKUJX8KC3/TBBOYNqWAhRysCjhriB720aNYUxO1q
H0W85CkOTIyIuB8mBmX4m9XPyHWoTj63T13MyD3EzEEI9mNFNDPV7ZhWLf6QOX4PRJ4MGcgeVNSh
3NVD1SWU25V1rLoQ2OtqLJuwAaWsl5t9Xjglc2IMlyxJ70GCy3rKxQ7dcrOjH8V0B5uLoxRTLDKt
+J0t2jfsEMKuyYyWiwF2kHoaVJYnmSNTwEooPLd+o9VWwMqhdQoRhp2Kfz+NCozNDV1UyV/tRYFd
3DpuYBPGkIIDEotEW6XeaV098h0ssIScfX5J1he3sF/tn0rlLA7MMMuALCfAMcx6c/cGRca3Kr/u
8yY4cGrOVH7XCn4lNmGxStAVutfV0xFHdySZ4E0y0bjN2EoZKpTHYeNAAIhIokwSSv6ZvUSej2vN
n3g+DVlFk84T8NxRsQIatLURSyUu4UbRlYiyaFOLEsSerf/vu6yPyhl80kJxIQ+4F9cQe82dceOC
e8w+AS/OQxGWaFug1QvrWPm6kKSq28kHSVeHqwKCv/tU4th12he8bNpGmxuNGsVMiDeXH2Ti2H6v
OIucqvGZk7rnZTVWjgDesRiLuLkz0tJX5/t9y8wVkKuFfb9l0ny+Dhng42gZ0D1aEqZwxPwh1/+0
9TxCrpzW2SqBD5gPHO1EshB9MtsBof6ngrhQfwxeWaVHH3e0yZb+rzeuJ3VCplIMP2MMqmk8HrTV
3n5OICw20R8EDKc0Sf5ad3kJnEvfSVCFLp+3O7a8rRVfw5xjvGkdywWUHxhFEIleJSnSEM6pM+3w
6BXH3b/teXXt8C8+WS76owe6P/oFl6TT+geS0ciH4wsZH45th/5XEv4eAX50wYcV3wsnYKKKKVOi
Tf7jA1pVBEg2eKUSz5nCXM/7cLJu0aSnVO77Ss4b6Sqk51HvJcSBwY34NPGd/9fKVa7HdiUr0tgd
qqoOo/GHbn6uON14HMkUYxgUcWOLi1RwmbxQlMbJ3ir3SGAX/iNEz1uilOg/EP6JDYJ6z/oQuwXy
GSLn62HYblIsfdLxTSzqnTgsRpb5LLuBeXv8lZIwvxtAEdoPjK969HqB3aL77lG7H4E4YuD6E1Jr
AhnNVkcHmpouvuxXeatfi1rsel1E/+9IUPpQCN9ng7XNtqemm341M7bAm4Vs7nNGMhFDtonvutWg
EY7waVxM+uZamDgDSePcMuVm+9D37g3ZZ0erQQjlhXZzWRo4UT9wGrKCLjdZRAjz1C6eKtbVevUN
42ao3s1wWCbwlsbkk4+Xdi7H0ND9Go7kwK1356KlMof6LS+CvvRWKsOdZABWIrHM296wMqDBEsqd
eoBFN3+pD0KtTK5DfVVrIiihnmwAdokk+HHOk+LAW+uEF/Sg7OTAdAW1HozkQ6XBEPAxnQ0Lvucu
EfWr1kqrHFf4HdvJ3b2japjP738CzLNDWMgFrQfei3NMfZq+cvkTn7vJSKtAWFG9j6+kVaZu2Pwq
2GTKGZxXgvEkKzVwEQdTA9HtGcH3nCyngm3iwWkL1BKoNBRhZD+0UkebnhuwNSzzIPTUMLz0gsx0
lJTm3/P8FjD8uBhFyo/PwDC1xKK/LFwY3g/Ra0DKzB1qa3gacM/8yIeOoEmtnMtoDZwqAl55mX4m
UmGztRJRNqeB03S/mhT3DLMQVZR5c0m6nmFVn78Kq/ZZwHyWMNhgFGR0ay0iNnZbo1JG/GrJWeZL
Sp2WYWPP7rVkeixBogrmAwo8wAp2BND7Y+wyGPWXU7ES4em8PLM5lNHcUAqYKqoGxg5O56qSYFPD
hShlul3AKk79MMw3j8vACAwDP8MMiACVCPjQVz9/10txN/YBeZDYWavzSmM09dux6nmrYkGTkatn
0FyccAM2NaTKRbigZfjUSxibToT2mceZ1ltXHOib9U1dAQarh1kQRHNcL/kzwEKLDsCB0w5rGRB0
ijvzhuo7Wblv8WjO1rXrjN8Ih5KFBEar+76hKVbj08Ka7GYWNdTOuTdy2XIvbAHYt7arrdiSvS55
bef/d6NS6/dChdIb6UMbWJA9ydhM7j8pK96PM2OVGAPGH9gyoF2EMgu025wQYvL5+AqXC1w++3pI
JvyMRsjQLvz/QQEjf3/Rh82TVeIjcibPE/aOIZltT87ooc5GKI8arrc8+q6SgsFIk20FEUsqbbqF
pP1AsNDzrBV6pGc2HdhnQExsXElk8iNUJ66kl9eQddsLUPeHzYmxBgHgGn2G4n1Bm1DceJ/u6BSM
dAvBG0CDP70LLG0d2w4ZmFjJ9f4C90WPuc7eG2TsvVgV6926kbI1A/crZUB0z9h4mq1OYeAReAsZ
wHW+3WvmHxgmqM9Akm7uohjyq/tqoiBpnZscq4iCU5dgZ14qf+T00ZE7acZ6funjwBEHvbdMYL4h
luSrr01+CX9VJ5ep5Ee+1k7vTGKKqD2peXNy8spwjTD8oCkrD5/uxWZ16DgRoBizEadEpiWcPcAF
yPkMEBB5yJ7lRgen0U44FPpAvcGPNVHdkuYGY8DcpOTvDvMtZavJ+D4/ZxS+zMJuiA1wRuW7JWF2
uCBqNjZuVk5hCwvpi10IQVxSceoYwRDFs3/pMSwOqsKFv5JlSm/56xmT+3FdcHfK0gXo99OgyMAS
W0WFVce7F+lt0/rsvDV8K9mhHaynomFufyrZatz8B6Jlhhfxsm3qblWhVJv3oc2h1yMJIgYi6JEN
9ef1Z80volS70TakyOz+Pnf7fqPJbBsV4RxoClWpOgFzIifwLkC1LfYcPz6QDO/fQWwP/pKKaS9+
lqMLT1tmmfGiXUp7yG5YwvuMaMvIvUe7N3JG10B/xpCtXs7m0mw4jR6cm9ZeJY5C69tqPuc92d/e
B67KEAL3AizOUo3fEvgQZLsgfP2qb6ORaow2cE7hbkonqBxQNtOZhf5dD973L8hbZ3FfcEjbQMmB
+azsnCv5+kgWi6xmU3+aIQq80HWiYl7bxaddzAGalZU+h9T6XZzSZK1hhIns458n5PduQV/aeZKC
TK9Z957MFvx1gX37xbcB3zMjBcY1qHHwsed6QkOOc6KWTvFEp85YvuLu91L9PX2xX8TsBJgiG1Dy
zrH0pdQmM2xa9VcaVC3KFEkyRv6vJ9icGhVHvbX9j7CWc2Yjd7pvffWt9zfi5AEOyLmMS2+yxPKe
Bd2y9FwUtcvcvUHp5nnu5Tbxqbu9HuWhesd05Fe8bi/FSYj4nCBCdy+KGqH6xxs4k8XRe/5q13aL
qEivQh8zuRDvqD2TkAIWwVMQ8svOLfOO3Ny2qzR/28fsBd6IDaDG/0GHXbHOUV3hNp35qPfrZSVu
rvYScJaSnntwvEXaL2c4QyQsdFgk7sCmbA0rwZUSGd7To7r9YxqA8C8f8i3TMMzimM1JsYXUejcZ
xvjOh1LDBt5B0V+V0eTKq9OZf1bSVU9bHTMp4+AdWrT/2qNbaNRgWejkCwe1W+VlY8Otq930enVl
FNO3nMNnAQ4Vr2aFhOgHrM/61q/aqdGGzLM9nS26yL6uU6dJWl3M8rzr94Xx60TrjzkBdZFSSHs4
Q4sgd6IinF4SeguFKSaSG5eB2prMI2UfW7rvWhbfwntfps2hi4nlIADb52J/TnmVFSMcKNGd1S8E
kP/V16G1EElsYy0t3rGj/CQn7E2v654XTXk0bwFvn3Cw+K69sEM3kqz3pmk2hoAw6IUFBmrUmjLl
bUjOLyDjBa4JVDVUveibrNWrjAtTvb+ag8XbrvdWRn3+tDgvnB99Oi3dgreswTKgc+U+gXiGdhAN
4sbAPEfkHzfPJGLaPDYNhV1Cs9JFY/i8iY8Malm6aul+Hl9fpYlktZ+rXoe9U7128X48li2rthfX
F3zhrcIZbTlQfAFiopxeFmQleYdtaaYHE+QByXItI+gYNHnOBRTskSAG3VwOHNx46suQAFKaCcL+
cVvLDD1sWGYR12QBi3MavIpyrDLvSjhTunnm5MnrArfultKnWpuYLJeAxGrKdzOS8BselR6Gy1mE
6Whx/CeXQBA48wqya0SfHbTde9ca5Ng0lYIvMN4kGiw1ah5FPxNIV2O2AiWDmJS+2X0IvC/DtRuu
dIsVTk7ZPv/MTj3TqtyrCEW3zrYmq1V4xaLLIqnTPYNJmY7PdR1X4ABPRJp2xLZgs8H8elvw1vnG
Gfvbam50Z1U/s3vrU728DBwqekjD8ilLddyvos+LVJmp1RDIyCVeBKgts/+GrrWJt5tf/WgSkngU
ey9/tf87I7TuRhUtGsQScZUWNCAO2KV/LBT+iHShJO4dgqfrhfZxTnDTcoNi2D804kSxAvPcNJsW
qljs4auAr3VlmkLzXM1uFejH2j07PbqS9087Ys9p2ua3s90HCMA5kUdu/qn/r9u3q3YIqwfMpxKs
WSG6b8mpJ7HHRTpb4SK8sB/sm2L+wmb4BVzlNVMFZGDra4m3JL8Vy+mrNZhgaymH7pj0lBUM/bX/
BVN3ymGHqaNIvuVc3zG+1fXhhQZrnlQEKXogFBuQxLM/tJGeN8wceNzrTol7/BbdvL/VJ/ayT4W9
OvPfTZdnblQAqqmvO4sbmj2V8HXMJWc7dOzZLenePV8tMI7aCM+rM1Zi+8drUOmcczmZywWlpsCx
4gEBj+3zn45v0WUKEfIrzK6U/z0KWkT3PMUx3B/SDUbeHt7y5I0km5AWiFZ5JoHL6p1UZjV0BAlk
v1iSqn1y3ey79CRU15Himy0dW9SrQ8/BZnOxyA1q1nwPQT80dS+tSjcZx2tKVDdqRUz2tC/3tJfg
keseAOIvvATncGSURtV972QFVL/ogPh07zHg65GBkUaWvxPZy+kRegMlXvzrh4McnddBJhjd7LIs
738K+X5Nx9y6W2pMXBiP7CZ2S1t8UBmVNzCk6Dw2c5k4otWQkCqwi2Tq6kR9JeaHerYOoEytOiB4
93mklkO3DZVWg32RTbxO4ULvMsXZX+b9S+pV9LuZSCmpAJ3tAY9tKC6wXsAO6wJM6l2YT6y9bJ6R
MAdsImoWnLuu+HwJrJA94u7b3Qt6mdXEoIH3Wj4MdJIBA9UK/mbVxGIlVSO40+USHg0n8aSzC+eQ
BtT48tNFJtQmUa/spIQlnuj4qt1+m8SOJioKjn81CymlIZ77wH2BZlctPtp1ULryEzctSAeOUBnu
qiRFAFNfKVMS+AzIrPnoV/dqRp6F43T+ubpNFjL5p+LWMl03fg5E20KVZQr4vlxUDHHAEMXgYdiA
PEpM5nZWx1jWQs+3xQWY+Qvd3xTuikUplwz7g2ZPlM4zqkNw3h5vU/wdmFB4sxYszK8qC62eEsbh
4hUPp1/olGZxnhc6ou843F6HHWFBbrWVgeU/G0QPAfOnHZ29eT50+xKDIjAsmUZN73zQnE2LkzBY
5iEIDkw/xWABgkjW2d7puZXTvWfxVfgTuOl7Mb4VAx+uH4zuIzEurmirYUUOE6Ste0Th1CzoxMkK
mmbcL2EjRYf3xsbPA/kH1raijeUaOYhMjKLIuRXANx0XdLmjIMW52Avy+4D+XbiTWoLd+ODAtVM8
xXvZGD+bjGnVTldYgJdZABjJLz+3qxxc/5NoO8LgbaXdc51KxwGzf0BxieXHeqADxSF9JFhZjX93
Fqih1eGjOfsXbSElzJbyop2mgO7XKYoQUJ8wlJDKo3yCj/Wd6vl6DlW439EqGKaL+a/ebWm8GyAl
VDuq5/7UaNkntkMMAGY95h8JoRW4pwc7zRQ1AmILVbP5J8OrSfF04XAv5r0qEP7xY1YkPtqr06uj
uG7HCyyFMa7VC3jmMa+H9HZz8uEEkD7SxiOevELLoQ9ZmJDeIwA28ReRfOw8L+/4ZmDehRCosZ/r
PCTf8IuQLthCjUNYamlPS5+KAmWqPuRvH8QSH8DC0AN275wnVjQEcZP/TWVLaHUuqGk1EguR6E9s
IxHjVXt4J4FMENkuY5mMYpH1s3PcsCK8UgCYrXEv2FGujw07stJDoYLUvqQ+oaQUt3NpXyrmBRKK
LA969IBqgfrxdGiCpWZXze7WBXicO6ScV2VG/i5zA4ZEwaBPKXNi+vLmQipY9yFZ4ePkjIRkKoqU
RH0+BfkAHUrUIlsfASpKOjMldal4+mj2gUNQ2TENKwbnpE9fT821RFyq3/jQfTg0ZvEro8yb949t
NBAMb0wucHpEtQ57V27I1+Xu2O2MrciuNXX7KQFHZDHE1G25Y+f+du9lcwuZ4jUKU9bdHjkRxQuI
lOHxIjLXN3PnrMTlvvhhjSoCQxQSbaz37IdMODMl8JZ4A0KT6Lnuou14ZF9AnBsL3N7+MZg/ziqT
KBgEexQMmOsKpwVfD8aqhgnGMXvbRbNdTgESjhxNiMwYTjN7fRODQDn9tc5g59g8K5oaypiAL9Lr
otIjhVYh6AjRWHyxr6Mn6B3j0pR3/0VBVvJL8M32Rq2xRZWadHN5qUjjucb9HlvFMoOFkcrof1Ii
VxYXtxSwQ0nIUCU7XCmtYk9sQTzsquDlNd1VVMyrfCHJewOjJDyk/J5Q9oRlejGFc2aCTdLxceWK
A2Ow0or0ijgLYDAYOWtSTpSkaPFdZsvVLSW0MOEyWBtLe9JG0JovsJYc+QQhXLyRNd1f5QpAfy8Q
U7W067ChEUhr7RDzyi/FOxOLHMzchAuCm80EzVHfqHBITU+3eD72lKE6+33D4901BBRfjtrljAiu
dhk6kwi9Tumc+TSDYcUN11/Qyyi/An9u9Uw7Mv5S0+B/yZWn/9kJMUtrUoRLoZPDGVzQeddQ20u/
NzcIdRFbe8F87GmEcvLfBl/1c/QWkLEmJVhY96lDWpIDLhfde0i0KNIxEPg3dS2tHR13CC5qR0fy
f/Mkly6cGxQY+nPLZSMe6r6ZNuj+Dfu0yKN/+PozUQJ3w5YHDE8AJjeVbZ23Ol4lIMWbe5gJGGsi
Yu07xgHwUnHMGTLa39azUZrscFHXcYe7qlRJFVTEv/tdIGhY2sbZvgSW12yvJ3sT0U0MhSXVWu0E
dQzyHEqcjC1H2VaNpncPPV1gHumsvJd9ue4/YIioV9mUgiRwtyv8lTRaBDlBf4yB0EnYoaqtJRXi
5exSNL3tvFc0J2ov2emp21RS4w444LL0XOPW7KEjabpc+9iSTZxal+JhWoyyrmsXQtNYxLMtxW4j
eQwAUrZWvbA/uDW0QvpDnirSCPTBJW+Io8lMxOpknpESsgTPl9PmSOMv6mcGrCwOwFoexwqRv0Qj
jO2JZi896k1oz0vV/8zKcjKXNt7yhgF5Y3VEE8TiaECxH8wUfN5HzyqFLxJKfoAnQzy4VGBB/n/w
YuWPxsr9872BqDbMhsoQ+SlRTyZVKpte5eM2tvdb7QDkXc7zdyaY6gyG/VXsa3MU5kgnHJ0Ri9yr
xDOPDshPcFZVIcKXTlLttabavab/i1yG9Vo4OejxdMBvAh7DtJmZJIS0RcwKiTRQc6ocTEpcZhaU
p1n+VraCFRL868eIwhE8WuZ8D571o6V6JZCElA/Jub4oYVhlI/wQDFKa6N3Z3h2v4zpYRnlQ8aU+
XsLOnAOl7X0d4DLgcPAaXDGnt/fEgZDSYhwFwzwhxufzboODjVow8QMddTa8KK7nfl36njaks5BY
/wtgHTHIwS4gZFkraSNi+AvYu4NM6gkax/0dQ5umMotBmArq2G0q70Kx0/p8c+LY8Y7O8Px39R+Z
0D9lTm9JVnuW4Svn5ZM76PaEmQyTH3puwBAy+IJ/BryUBGO0/UaLZ7X+6a5ED7llAS3Qvhx1Sj+S
5ASg5f6t9Jb7P4klRQWWjuxuOFXxwIhmSlXhc3AhJF+aDOTjxSC9H1EldoUNaceCzMBZ4YPXdASv
119xI6/NNBxo2i604GX3tBfueYeaqSJRxeyQfwybqpWJiyWMHz+L8kf32/eeOR3i0q81F8zOKQci
DjmIO4EiwTLuCP4XKgnJtRbwq/nMc7xZa/Eaf/lQY7kznk3WdyiOGwPpPPZOKtww391exr1gtOnc
O19VBF1k+0UdhSDhOmNZlU1euS2wLZ5GW1gIyUljQMU/ineScBO5Q/4hPYsussR66ejzmwVZzVLe
av92khocwJCJc3ULvdvmDLufbbtloiBQO/yFgwZdSAhqj/zQ3gDMtUIQwP6Glm1+WDlfVRu7lx1Q
r5mEQHK3t9aeBEpSKsohuZCTrSfeA9mR2X/G43MFdE+iTSieRnVlTN/oPRUDvuvxNNbBuOcNLR48
7tDXo3Ma4J1QXHD3dhS8kp2nPv8Ijjm6JJIKhGYwNX9Z8S489Y1FV2HwWE0zwgQOr41MEUDlNDD3
rCiLIsqbEbX3ddTXjtAURO2NM7l0j30hnLwpvYNPZO7UyDT9AdL0p6GMpWYBgymsWbvGJFMIL8qw
3pwZFFgDBuUoD6GBkQVCCfy11V9ugOJoKonvbHO3QgRGmt/gndAU+xFVOAKfP56kAc5Yjh8z8TBR
Yvz3A4Ej2YGMrL5QRPoB7DJxWVf44SlPLdbQ1Olk1o9Cl/diurtubenVr0rwa4rdG2lwmGd4+N5a
0fhSuUWGL2ckW05M26+fOGh+GMk0sfbv79sswdwkZU2K+MOicG662w0UOsIyOz34vikyYy1UUU72
uzXjM855Q5vuy3MI+z8HRx0HmwUYZzmjDqBiV2FgHhqJhcHWdN2+P986tmWJsmfw5vfdQU2pJoHz
oCCuIxlbiySMOyfaK5h8bER49GhMcTHxeo8S4I29Po9cGeEuAGIS79HJ94h+If52jGMgylY0fsi4
SfsirisrOIqRbs4TeQim86srsCJVf8YzRRrESI8VIqKM+iyuA/QrAaOcisTtMV0kjkJfkVtXI7hM
iNGG5/Ni4DyRwpOr7kZgw3bViAkrjJhuArCemCN3e3iWsFq48j7Iz7c9hVY7ldDm7CN7mZYbz+sY
ExQYS96BFtpQJUQ8+Jk+JS1vCSHGWAq7UNglRnc25LKJeMlw/gAAbv7BjxJCJ1+N+YvnmBvaXK15
wtdPOHHBMAWwvvFV9JUTOa22UNFdjGtmJFMdwG7An40W8fxqCJ7SrqxkRQ5f5fV6WVkIsg0VqnOe
aG0lXBZv2ULUlORvtsJH/tYvqMO1pt4YpzFbTbmM6UQEnUB9LaIqn2moBJTQhkQ3XygUU2QI7MQJ
oGVINZsKrVZEaTwYfIlbDd2iAvGyJUUfRjKOsvekLUM1GlKKzUcVDwtHaKmeoMTq13nPmvAVzOUp
uv56SMf5M+8AcQybv6G796D/xY+BrF4Pqy7c0r5EeWEDCz3Kyhs1gfCN7PXgwJq9E3lDKfquACwE
yErehybARltKQrcgZGI+g/4l5v8kuThi4jGQ3deebZM9UOQypVgMo1wgd+DWKL1IBD4bHhzsZpro
JRRilJybUMy+eghBeVCHPbTKadzjqYkgP2XM7/m4JTTrthojFqIoLIAaFZUd5bxUj8f/hgqzgksS
UZSYIBJVXsbiB2NAd8b99srl29961nRr+F1KEo7lEgr2C6VeD0q7kVu4P/mhUq5mZwDWN4hLE7Lu
SnP/Wtu02pfZGkxlv8H4K5g2Gd9+gry+NQuoIxmux7EC/yFXf25xdHt39qRnDH4PYukIdwZdDu0W
90dN0dpxu+5BEMqHiDVCEKnTqDV2a0O0FLcKTIue46fiLbr2AV3RhMsfmzJFmq+yIFT4cddEdHwJ
IzXHg7ZwMJJ/uDakrPh1ymFFNXUf99pG1vn9SJa6gGfvYF/Glajrrzb+IHOY10n1xW2vqSJatjpO
j8HV7NxcwoilPQuOwE2WG4iV/p5/u2MsRAYNWf9WqHadwjSc3YqiHPOh1aog5t3rk2k8jB+8DCOO
0mOni2n7DaKxeTYg9dTySKlthIzFr6R1WhgS6LB891uflLWk0lwCvxneF0YyN8cuRg6mzU53y7nH
YiqyOOaHO+XHqV0VL1AMKGCFX4+Q4VudyYXQnEx1QJtfzZ08pEolkliSROU1VWdH9SgGBwu1XgYw
1T7Brk1oiHdfcXTq0DdpCJ8SydESrlxeC1OdKbF9kKIFLqjfkHazZ0P0k48vSi9ffdD4bU+Oab6s
JauxwRfhVo525QdS2vigVj21v2cwSSt/JhBNklSw1SCtNlgoVAcxdX17ZycOSYdFR3mc5rQRLpJ4
Q/WD+dSmdlVAXZbYLc0/BeW0DAHEo/FdfRBQxUUwf8uSMmXe+Y9GTYzsCLXcJXZ34jUU+NOaQ2mD
UidvYI6NlKLKBlRXlFyG/l9WRTBMISUvrpg+PKLUMEzjMyPV0W3az5vjnfinukcHbuYO1hBuRJQq
+30SVqXKj43tYfv5YOQV6i5LM6Egd1D6qfNj3r+aMN2XD5x0BnjeOSHBCAoUddFya+yCI6nwiSD/
hhL+cFk7ux7bvXdrxlGr5lgNantO+DlSpiiScfW6sgbfBFZ0BrRWtNZ28pUNJeAcWMLS/fCHim8i
IfYAMcmSxV5e8l51H9Lw7YXpWGuiXXid9V3/c+yoeQ/YJtqxfUuAzbgB+aD3RA9CvxENrk9fUTGk
q8tS3eZlXUAkuGcO36uykAncsgFJrOjsg6s4/2YkFpBFgAohT251Qwft7VR5akukL0wGRfdokrA9
QdjLQFztJUw7MUPpdgFXb1lZjx2pJflG2fKNVponKJXQ8Q/pxHUUKPs+L8WkGV25itPsP9PVLAhB
Trk4Hlln8C68dPiLD+e5aot8YJu0EbQkfcz1U0KAbIJu8iomKPr7cxxPQQ6Q/ZrULT+P1YdQahs/
3pBlVVnRabZi8B9fSJcbWbfgnlhtvrZnvpsIadFoUCIontAtr1QSXqyQUPOyiQ3IB8c+sfti+d1M
6QjXmdCmOXmpoSCE3qVUGJ82xNNJz+JhCgea5XWf2Dhd1aIZAg72g5DJcurqRQG0eRAbrRSCPSyA
lCHTAh26pLAtroAMpFgkRr57vSQ2UwkRS+NiFIMJqrXudvdF/HP+ytkWlTSm6IScznPPbD3davxe
Y4yC3XC9buK2+j8tXMxFczxet/DeN44IqJlb0X6cx4wYQffHiTKgIeEGob9rPZspZgezeSQ3tQD+
hqCJeqQXNFVwra1JY8UB78cqErgobnkzge3gbis5/oRzmaTfM7ST5PZohAupyjd2Kt8apgokH5de
YCFxx8E63myG8W/6UxyNc9nfjetpUhTWHM+R34E3DfoqVUXtUq7wcQBPAcndf5jIF+uTQnXxcitB
uOpN3XNtV+KS9VSzvYyUTUNKKPItTM9N1j5ymXhLQERofBBdf2Yoz4WkbfgfVYdQ2kmANfH1usTh
i7adA1J4D7dt3Qgqd8pmWW9LXGJo4abGSDMJBgseXjpEInXuafRGjsUvtHn9ctKQkyfSMfyuK65o
ZeIjJKZ+LRqZxARmxs+PGw1V7WqJ/1JoqixdVFiI/xIe5dojXIwYKfq3ECXDfclAqMJn11TMfumw
CPXR80AXfOe1OPo0BFPYU4orTVTkB+96uYcN6zHX19h5lc55/PckDJFtZa3CVCsc0IttNaTOCuZ0
pP1+Fq2z9B9To3HpRmLTI9/Rj9gVPIDjc4zISmny2hO785ZWLNM/igkJxenQr4MQn1JMVCkqmIlG
OE+AS0mJGwVSds7F0KtQVc/LxGMvsZHxJURStrqMDvp2EU4R8tdPi/IdxZF1jRjwMCCp3rMQoVgJ
CGYGUvX8b6FklItquPzPWTrnCPpIYLiVxOqhmkaHjmeSvCDNWHGv4rIMhdFP99KGII4PMY/0gSAu
sb4HcHet9PHgOrvcwCfXY1gfws28x1M719ETjK/ZNdtPrvpV1WBaJm5yQ+xjyigDskkG+I0rN+ct
s3smcd/Lg7fnFDkIUof3R7lj7NyaCSj1OnYnp3tSfZ01jdoHY402Ave5qzQREcngWUUsWUpuzTgr
DiDFUDoNVZzaP+1yAXw3qdZeWl+AuWReelQv8RjikSSsaUrP4rqmDbHn8WiQf/6Q3VwxY3wNae7G
Nzi3Kz+RnUZZpz7rkXFWtpFs8+55hbGbIkknifj3QizpHLbKnHzp1IazIss3N/e6FblRePYRdYzq
n9tgEmzCEvzvIWeLyfAGrq0lxJQB9ct5IJS5uCSnldyFqj8a4azQ5NYEYn3kqt2pioKc7YTGZCKQ
M3JUkanrNtn2WhEtylGlElwRn3ZVzjK8AlxplwwTrQqTBf7Evl57ZtkIJW7L4xxO62BCsmcYANH1
EX5bi+jIY/qXCi/e0fT3hm8Fu5jAtzhnGWyCi/LUgGA4qfXYf+LHNgw+u8eO4jaPRklnw4lzi4SX
lvCCtd2LKgWygv/KWVb9E2NvNrhHp0WtQ3CMcYPAsoo1TWSy+Ui9AP0e6grFJK+pb3atpukMH5aT
QejMm6NNHg0ZcNCqku9ETDk2SARi+6/MgmVELvnVbQ3ySLZww5G875EaVymoMTqnD/ualNh80gCB
ltwLmtm3zdEpE+0qPP8TzM/o+tDe28Tl1cSKdrgkU/fyotnd7JuNtPl5TAnAoNuizKXnSLHvEhRw
SzWT/R3ndoW192TygG8jBkDsm/P7Imh7Lam0Fw9QMwLW026+IeBNIp3gSjThDKEFZs7RRBxN2aHn
BgDPsC8RrLnmhIHCZ7BwMPv0XqHp/+rk7jQuhUiNSsLJ5Y/emIWQ1nhXlHyambRtj+a1EXDuIKWm
BpXl/VL0cl8i6oYr54URpRI6Jnhyj5+rW2oFl80Cyr6F7HQT0XOvwfERrvRTULdaqoF5a8d965S7
6c8fIs+PyBsPzdOXsLpxg4+OpQRd+T6mH8H9h3EYruFQPvwCYqp9iY/Ug3Ivi1B+LiG3GMdd8E53
GyTQ5kXpTx8BB5jxLkPanYM0cUFBbJFddK6t+f9fmH6rfyTU5h+rvSXeEbzcM4jkywuwSGJA9zrX
sdA7IImqkorFlYVRPWdbyxG26urpwPWn9vZjBp8ZPHKYkSB/rwm1cVBJMUGsDX0JNhUpnV5wMSjt
IItt98KSyvXM6kViRji3lJAPIWN4a1tAh9kL1ybJrRsgFMIhd/XnazZHv6L+iBBqLWcgMx9zYd+9
J8/NvGPc60M92nAZEqOvxeeZnCUwHNGDMKOFyn15v0+jVW//Ae1shjRMjYcelM/ODHLkmBx0QZpc
d0LZjZXtFp0cWEQLb8Y1qv9BR1higu/LfMuuLnH5CjKnraq3W5hBY9BDMX10FpJChMKhe/vHPNNV
L1Td4BrOCSOoqVTAn5eIXuwxwcGsgS7Gp2bKJ5faIGW8HRZtNqRmTFGyGBxZy1cYTrF7ZrdqEN0l
e8VVfCDVYr8uNwB/oxY3FOdZ/wxbL8vatFt8ctb0Gg6u9jKJw1p56xdT765V/Q+wBmADJjj3mrlJ
EvjFRWIbX+XJzplxtFy8pQIO6uDVqmCm+Ni07bwaI4VCOGkcErP2k3DouG8JrrI+mkL3iNIdbIGo
X1xwI7NC+1crIg4ArdOJsS5WPQlWpSyDc0lk8Ho42txvOSSDUOIDL0YXQpGyX/k/EAwOIg1z+HUa
SRYytnHIBkeymyUXIBULI5hQvgcIT2DSX4jZUngRvHsyy6XbKgPx6vBx6E2rZzhidEFo6aZKwRtu
W45gfgRoaODQmnJv7OOGbFA1GldR0ESHGqqRDfTN2DUjNR6QXA7O08oyio6wphPAv1jauuJ2DmML
2rOS1chIQc58iKwPH7hLj+aS8lG4aBfLTQKWLfUO3gQZcI2FK91VcYb7zSEaqkE/LoQ2Qj61w7fG
jNZj7hKQN+eF0uPFR0QA9hVnrPzMouE7CdTj6JGj5kXdoUYpYh8UPouO5ApsoZ0jZgb70kFhHHc9
o1kAIm5H4ehm08ZPM2Cpki0dk/2SaHEsFeNOGdqja0mViztWb25cWXAIuE9dpKAtsuoRQoP0Wa/Q
WZZJVyShvdA4ejabxPxTcX7QQnTBpdkNuHFlRTpST7v7ZZBjcWsBX9FrA22bOtu+i7/cmQYGgXSG
YgYGoVbDRXB5KnvjV91EseL2SI7L43krftg556SlcymX1qNpj8kxoNBfpw/Me6JnwfXv/5OHeibi
tRAa5aww4Iu/U6V7MV1VgfQrf5hEZlJutpZRr23bUh4G4VM75f7Ww/VWDcEzM6pE3AAAHjzWtlbt
F6FzJ1XzXPLyfZIo8KsW4sjWqt3nG9ZadTnkPwCyhifL+Wvh/alHERbJ3RxGuJEY/bL7et54TTs9
wiomU2N6AyNmnhzfwWk4KvD2DPVXE/vrW7WJ+lhVEVixJnYcOmvTgD6oxOduRol7dHDK+KLpR0dl
1KXGw6NDByCDUnHK022Mzd4fU6deug7b8M4pPgpBGqYy/3J+9uafW2xu5MTJnIExXjgNZyq5eJHX
lGflcXGqJv2YJyvNXYRjlmtIuRwpxgr3fwPF5sUdurpRRKsgkLRkr7Aa4fVVCj//NFCvgsvAaKd8
vIo3W6Aaq5TpXnVsiq2QyKxH0JWyfv9BkHf9AOK4n11sFKbFfLYNTtHLGUJHyUIO6rdArjiFNmYc
AOQnHJ15tk74tPVFbI5OXyXHH5ULVSsMk8WztRk8knazi1/ULhjxkX0MtvuqpzZ+BqOR6ejM/N1T
iOQI2Mxv/Ncyb6TKP5AzdCHgmEAWMB2GuHK1J5Wc0WJ4xeZvkWazzH96VAww1JIwjr4QUgfMEzSL
jrz5guiJhL3+66J0jnhDu2PP2MHxY13TWEkUUgSOLwyf1C0pZKDFmSWZlB53HFbARkcxxG2IkYvJ
Cxl17V9JRcDokkTtb5km0wEmZxqFRfNsJnqUuXpTOjmSi20nJzFLAK6E4ClhEfpf6ZKS51w1xr61
cYKa24LFiBftJv//5Dui6Pwif8lGSZqsM45+FzYLQOOLvsLBjA4i6Q8TMGZV0qEAiWUv6W9JpxAf
AqxnX54m7uSuDLmEJL6Lbqh+CqDewGgY8NJ2DWz/+UIDZL2EnbIk4hl6wzFnlf7hNZeZj3DJlSfH
K1z1sy/GkOu91wrGNJLkMfLWf8+k3j0vY7runSnC2SS+cvr4DTaqCT6TLj7xTktAbqC0Ofyc48TQ
0gH8pbfq5E5vOosOqg+0FEA6ZbopgUQlXyGO6HgDijfvwRi5GSRbE36Iw1LKFI9HBLi9+nkmO6DB
UU4hP39BJcRuiXT/LKJWhnFzNEryZDm1MkRKnNgdEQvIJ8gtEo3FJT80i0MjN13UUHsfBg5Ss4lV
PXQ5QggGPl04y6rFM8AAmayocuiE1+aHTahj1a338jf/+yVCO5ntCiXRTLrtRqUolzw9IbSc6tKK
+Q/yPFIIow7ODHz4cRR1oSqtVIKBWQK3MdL5ULSZgMTHFCORZ7XF4A9meacINPwl1Y281EOoBogK
rnbmnhzL3sMOqfvK2fHBWMIpOg42/aVtXhigZxcoVbErwMYw6yn3dlpxiUh4+1ZF7dAC8gxqxQQm
NZtx6NfmXnW5d728C3WeHsJa33YhHtQSPOLa5OpH0muhxxKx27zSPY92yH2mmdwfU27iAFGrV5+A
RZSVfYRy2GyVK3uCfnAEVv9nWaEVuZwEwvBkTxdpVsqzyI2zrxwS8uYKlehmyoU4AQ9j2DH6Atvs
S3pLkU84JwhHithZiiPNKaBQFwSef3GCAQSFomSmpI/tRGoHNVxkvMDFr/BvTyfxRMTOISDSXgA9
mUWQ6huhY/2W3GuMcoUamjIRpD1EExDE4qTZuBqrQQhhcMixvn8GAilNoE8Y953Kpp8Ja/93Qjsn
7uVL9N3Ngcd/Dqx9mKiEjlKxcWfFTTIRvJIu43ziSy7RTx1UqY2bGYITdFZ5Oh5C2G5l8sda1Wuo
RS8uxT1djQqVKJLttyFMpiodR734bp06fJq7EuJJgEMTV1EftKwmQVINzNRWGGHygR1BflczodKQ
eq4o/QIUVXYsFhOOOpS8/nSj6PEVXidguzopsYoi2pELciJi1Hnayv9yla6Xhs39E2/UXIP9wRNa
viVN41XTzauNGp+WqucSSi5u0MHzEs0cns3euji3HdVeMoUn/ernAzsOqK6+QfUdANjFYnGlZr6/
DXJf2npPYiK9bSLWaTysZdNTQM9oPpyg98PNeH6XgYDX2656f9Z++ZvWLRaQdJslk6XkXHiT8ZYW
Dns8+ft4gb5YHnShi/H5AhLUU9KsJCmyPpezgX4yqIaOloQqO6L7WhkjZR2f9hv3P9+iFic7LbxL
IVaVJERyLmlF9bUuHCioCpK9Hc5MW1bHe3T44KMi5xnk2PH9k4q9nCWJtZ7tRqe2O28jt7+P6a6F
Ald3jXpfryno5WgdLLdmwi5gsdmzlUdBtl8WZUejf4FqDyQpKGUkrlp9IWL8FzqV+HaC58To7KNN
8cgvSFKT3LrhuMsEBCBpAFUG0fTeYcN/6ltq+3U0Xmd8W7PgJQ2z0/gAuIbg1n9aXIPsB5UPoxtX
5xxAaApg5FZ0PIlPdFYyG5Ls5+CSdxwAoZg6yPtn98d4u5+kH84dN5/nIKHkzRPZKFpYM8yhd9ex
BEPt1h99ngBmi4NwTRXPZAZZDUpQSV0yJm539CPbShhSra9nMG/KZhddtvEsN8UNnskvkSXi/H5n
HFLRNyKAZMJkt/eVpKcTb6Gqg1sX3H4NBNoC2zerehJ8Hvd9NMcfGFAXTeaNCUvaMnXL6lIUb3Gz
f+4H+ad23oEF/ZffSmwMWwP0D9Q51Lq90pYSVUwhdT+bt5wVreVTQLFh99tOIdBNphZUp6hg9WEa
82iERucf05S86OVvwhIT/QfFr0tbeBy1Auw3B+US81lKgyfWUJ+DXvc3J1L465Q67jdiEyhuWriT
lF/fombNCXjsgxQfHONbdlZ2aT2RpVJE+jmEcQFVFHwiWViqu8tOT0/X34ob3rvuNvZm89QUE/aV
ktchgcUs8xbcgnSung6RAJzFHwKGNUkLwkC/0u/1MLuSv9uBQjeIZUpL2ZDdICvEbSQAoEYTuh4a
Ttpk4gF4fgNpZttsKQdCvXY0YHOk5Zf20zBseSrDCnP2xH0bCug0bYpIHuDGUtniNzX2dnQqEFX8
SxT9YowWkQwzAAlVW079XUdRl1sw9b0UCupCYm+GX+4kqiObuvw+usVMOE+MYs//iFbJ6of8535p
vlaPil8OQriHPgheb0tY8GDJT2natJPJ8hNdgfAC0j84ps/x69S/ClRo1WID2sW9E98JYMqRFC5o
9icP2h+4Eyyri4JUBUR7BHMXTO/65F72/Ix7Le0Cq4JFAtL7sCeTXFTKotna25+5irGnIArdEJgs
NhmlywUTBSCDT1W46YWneHL5XK7VUgkqga0yitZvoVwvRZkDcphv8lPOTnCi3mHUVDgzRLipqD6P
Cod5AbC7FufmbDcX4tLs4NSnPOulq2IINtfrCXRIl1y9zDe1kNMPDb4zth29dbuJl+eyXYMZ7vNY
X2YCn3b4f+zaPLTSErQtnTQVH7Yud+MuCjEQsRj9W8I98+6JETVkcw/PQ8hSD52Ht/RfIt8eLEWG
6xQj2SCH5mHZG/+e2blCnX4RBnHTkW3TmRTpXkz3ImndHlyUN1DvLqbh9pIkvOtaQSVrybLauTqN
wxbVpkcck87fz1ADpR52htZxcA9f+uUyl5uKZgSWmez3ib7CKHRnYM55rFBiQu2ZqCU0zm0alu6Q
VxHal5G+50kjhGub/LnEZOeUxYUOKtZzf/06KCgFpAr/ZDADx2iz4RVZJwebJZhPMxTVkapt+QsQ
yEedrqaopk+75Gvwd+kDHkOWaxpA6VFbU8sPi6is6HZQa6xN0PgCiqmRkTamrUHMaSf2MTH6JReH
U0ga6G5NT2t+t9MXQwdxwW8qIcXzawfWiNTi4rF2TkZmqO0sc3xAd8zH/lgpWLxRx/2f8hozHJqU
NGCR2uVMTx8VvmO8mo4mG34M99lATTfZItEazg7o9MF0KFc76xWXRS8S1Gs6l5loVCTf9fBN8Ufm
uQ93O+Le+Q9q8Phj7/mcSADk1TQzIBmtnvjAXOmNqlVR2oH23Ao2KjoI11WIj6AfASiUtS1bB5SQ
uBI675tshoT7TuhhCqWuHNKIoCyphT/tRfosvZ8A10v2H35HROuEE+Hy1AOLC1oo6OIAKMUW/4CK
fI4G6C6MAlpon/4x0/Hi+W4oKE4DUGhK/Glq3OMj1USd6hvDwcBq3agpUsfcXyozBHJq82Apjz2J
4ljPtl6njFYv2PIyNc7WLO2OhNSiXXi9INkdgRSwNVRzYWga3PQih0FvX7c9oSk6+DeiymbWZSfF
ntX5xtT385V4Q/Cpsba67Z0EbrSsawfjb3PK3E++qerF7aR/2bCG/YDvaoEOOVNui/Qbv+hM5hfc
1Ubhox9CW22HA2qy9d3BFjsxQ4gkH+j6bgRVjjBnMKiwEDiN+HLqXa20ZxBIdgfg9EWHbucbti/r
r+aug3x5EDTdtjdz4zugXwycFerXTT8tR+Ud+57DxxG84QsGGtrMxpcHCF9Yv7LFYN/vyhR2/Y+A
Dx4jMlBMEfFrsXKvZQQB1T47qdCORmRyDnYbOQIF9CiPGjWUw7JOClKKx7xLllDYMVRKFgMBQM9g
d5/puTL1sU4Q0WNl47DhW3qLhgjBJiGnqWg5HdRe+2n+CzX7/1/xnLKIQh5CFOgy51DHCxank0NT
Wrlze4xhxts+6pDG/No2+aHhU3QJg8fwWY9585faksdAyIj1hOd3OUFY7MkOlg9I6ysycA1M+cgm
VRAOtC8nhtV43KPLZKHOjT+yE/r7/yhqtKNLIwguvV1YuvdFAmdHu9gG81uMFRSzkqUyX6PD9xzf
seyA/ybj10JkIKOD0GNwN5iFCrBEjyMI8Hirw345k0d6CVZqeA2JCZfyXPpsisVxaG2enWHB1gsY
jQgV9+5s1YFvf6cNQOcfLzQYA1nyNp48P5a/B/cn9PLXqt0cmSU6rkk1Bh0Fc0ggBGn2O02geO/8
bhttKwdqlnXb8Cl1/TgljxVs9tULNBquYYnT/wssdbdleanpMrqDe4+Otz+bN9lwipN8t399cLV9
sIXUGyrraKBVjDgjFFhrK1RqRwY2PSggD5YySvmIBfAKwz2X1vN/2aFxRAJ1XPprxBOjTjwNdWO7
BpLnTAeEWGLFpVHXB6hS68NMKoMv8ZXAqNidhwYLqwc4AcCMAd8Wh5NCfhNNzw3XP9PFSvbpfbW9
M7/qbzq7uKlYg+RC09/8nw2eW3/CBOCA2WFTj0bB4j+4+LqCQ8iDJiRpRO9jTorPrIzGLwtVQLxl
DQP3W7+kyxVPnlD8XOSVtBk/VqnS4ouN1u95SXIBpr7bqhMMBxWcHYcTHWVTYT5NLJZHsmgeun0D
LX0Q3tBRZH5zSGyUr7KW0oE2cv5KTG9TYXXpoml+NJCvoLEmq+48+K5oYltRHuSwsgkrvMrCQkLr
KcGPfrKEWZdyFE7m3854Nt35TSFE/fonuVqeDaO4DbFCE5sdL2rne6JdIfsZwXcpFNu1PvdIpHhF
UwGs/a4SlF2QovbL3tJDKfA8haVVEh5sD9Ypi3SKi1aHPn2IznGKd1xr7CwK5DIvEQbdeiSLYngi
59abzTh0hG4j2lVfKOLsDrbzAhkwTlZzP6rWsxeH4OMtaNdb9pz12ypH6txNQjm6nHddafW3C9k5
5IDC3u1KNebyQo43Bp8ZN5P4+wLAy7P/hIBfq3CpqllSIeBPxxdJox4sDeLD5nlK4oEmkdECA1sZ
y+/phr2BLJKUdYZqii82yRimJ8yRzhXn130HZKEXEylr6oNsUL8J6wPsW4T5+1dDJOlBQpiDneZU
V8TVG0qx9CPTqjX9Ltji/rHcwNtYQdmdML7a2xErbOy0w7kEzrVMYkE4THpLESLtR8MKMW4Be2hV
uH4c4NLgDEmBnkA5I5ppdq6KbvmkiwzCcQJUzIFJlx0wz+N58OKJPBwInDLVMfZt/yvrK3is/KHL
ZtLEHcJmzHreSP+h0G5PnqWA7zLNETgbQL4CEeVDJkEb84wTJohN8FVDHDZ5bMpeGiiFznxDuWH/
Vnj3jeUzIgVpLrKdwlX+StxcwFpOtmyXMxeHoJdfL1g+JrPZKDjsa92mzyj+gkdRiuCZEpoehpd7
hos0mskyiuFiwloNtt0XoBvkpFokrOvzXCzw1aEDaM2pi2YqNnob8aKMMky4X0wN9h7JeqAUrCPh
lzF4q2paRHT8JABaVI8qbv/AtaoAGMpS4uO7myjWLbvUQsIbksmmB/+kudI2v+6RfLr9oLMJ9Um9
4ft1Dm0hnNzdan6YGNxz1jl4dVObVHoUoAs6FTl6CzMH+8Lt5W0CJunXFYjrdqHYPg0d6fGKTfKr
pphtkeeSUkAuOD3bfIDRShPrK+FiIiLiDnxhXp4tp6X7Pp1Y29sQktFLAsJI12KOR171xvZ9hU6C
ahhuy1Uh5Ny+fKcAnPKK/gQSuzRnTgos7PPCKZZTzINT5t6UgBmU6uBw3cz72L1DCP/wFbz45yEx
q60AYL4ev9fZ79E3/grsVOPZZHgxX1nVsgD6+qVzOe/tytIQ7sKneatGpQj4u9iSIz3Zn9hl/5Kv
bmkU4zGU9xVZym4q90AS0ODnEcL5IdVlFe4HAhDt627OxYhVL8tZ7yrPLRZPy7QQR+nFg/TIr5SU
0w/FOQynNgz/qz8QujQ9HDNHptsok0SyoLurTGr/cg4QBq1fJZZzUw8To5eed3FzfYOpzPwwGSsI
qw9WlVfJukZZ5PcKq/x1TRQkrwSSOt3/Waz1DqapUgdiQG4282D4ZeksYgJYV00esSSYQnLSLv5H
mSjzztoKHKlDYaocsG8t9Q61lVQzxNmDocM4P5KWhi+cX/1ndvgPZJ6100kKhnlb12Mb8scn9mYC
duoT1KRwkXBXaqee4byB84jUZu63FJ4+s0i+Y1ETxUdKxa67B1c52VkGMPxvrM1+QV/BIT2410+s
w1SwfUWR5jpc45fSe/YDhV7fWS18cEnxLlb5YEDPn1/dAT8D17sB5hxOTsT/zPthIZwKrZlEBFMa
SQjLDvpK1Wak/+Kpeb5uKhImiCrv7iWKnW8uNAaI7ZIH8DFLwcrSohFx8MjGb1plorivqv7KUOt0
JKiXT5C5t6r9n7NlgkWkTppgrXtfdSBV/YGAfacKwvfsTBiGimE2CvqbPkBuhK0Q+oyTce/YvYBX
8nHfH6ObFdKV74OeAUVNBVkPOT9FFDDukIT8S/F7I7hkr1GX2OjZKdH7vRNzNeUOvhhRwxmrquMY
HHg3STVVr49V9WlJ5t7o/nSQZxDcwNLyPIi2lp2XZS1L54Wje9VwEtjLVNXrkdGy1Wyxz5WQLfIB
gMcwZgISPqxnFLZhFHEAgUXkhvt7BIFV866s6Vm/uculxCMAADUyolnrATO3REQrx4At773auUJa
Or39a7IeEuY5stmKgkeaI/kg3TbgZoAApBdXs00s3x2Yi/cMlnglRGXHSfbXWS4witRDF6KpnBNZ
jQqxFdDaTRS+zth/dYUVdubPsO4V0emVFVG1pYHdC3PuG6ZPg0IpK8VJhhyacMNquVOErAlHlKlV
Z+snz/CeLj6LT9c7VwkFkdZ+GlQ/SjkligE2v/XJv28tvIGV+C2Shf65c8r1PrKTmgLPxbsl0kmj
vR2UXZ5Q0bcUIt9a6b8vifLsoSe4o+zm7p4+effkUIZdKZojQ9aY1xp4BQZ/kXYoi4SGBNgpSaX0
zI/jUYp8SoxeRURGKrM6/LYZRMW0PD1EIW2P4vHMB5/BZJW3erhNwY0XTfMjMG08GS1o/IGZhrou
pja0XItACOb/Goq6k7ioG+LzLxO7+ItSpqniJH4n845Mxem8tFIo8kClRN8qor4pl0uDuywiXrfD
pJQHGwXBDL/MUxfnk2PnHagNCNJWCkFgnmi/wmmPLfGAmVt4nOVYeCIGOfqgOYYtasve189Bx9VM
vQ9tMxI9Mjs0gl6JghlMEOLytg0LYFmBwUPkJXLO+HzLDTC6wUc5/YH9v9FZlYmdbCecQ++pDOlT
mW/vzoC2MU0TY9gsz2SF86L+nffVhS+XwmsEaCH68yRqHHq6BMmriVZh/wyz2T8k18lxE1s/fQf6
Lheoi2MdKPQeadTZZA4r94la5aVXTK0gUZxYbzi3x0Fr85uB73r8F0oOOoriV7rYSuESihKvTOQF
YOd2EVcumCTV1Y1lBNBOLDoHwKYjC9DEE7y5L7FCjZ2fzyDWykCTtCyoMdWVEJTWTcHNr8lmeWie
xsrsittUvOsj4pAvVVMSeLvMaDy0ZiRJUqnusHM0SbuVqPawS0XMiK64MubeaZhlAgOAEnaTTMz+
meHQSXMo7ScZWH8nnZrNBaVqxWoZx1CGT+MAXu9rgu3GPpLE4YXEXQfzndkMPUuCW7NS1uXsbooC
S9+cvyZxv+VAs97rMwEpb8Oum/hUba93DC/HguSy7FywzROrc1qdeLJ/m0xn26gDRslgfKGcGGVl
0ePi3VeQgsHaOWvJI4fHlh3zyyxWAh6Mq4sjP8Bk9xPCu9+7XWH18Z6tVvbBGFlMRn3Om/YTDBMq
EJOKr6z4Y/Z06rl1ayg+IIYXDX3PFA9og+LPLCN5VrUm8A2BJj8EPbgz+QxZtYZL+AsWt/Dg2h6O
wRYHGLVZd5ttBMe5WeYK6SQeH9ThVtGpwDyZpqBkihc1kFR0PBTjY9dvkrovRj3/lw7UKLndlNb7
rkbM5A4bFyrOGAzVoTg+AbbUqHvNSv/OkYWY7xzo4qwkPlNUib0qCAg//m3xDpNY/KgClAbk+7jM
2Qzok97g9V3za/dTwXYGKIrr0Vq7jcS0sKKe0cVj7WIzWSHIOEN4Eb5ETa9a9tZ1ntPJhY3B405C
OmYcbzSd1MlXQkKwqHJu5UpYRd3uXfPgcQoPgw1kEX8SY+Ze0/5UdGibEcZK0H1et+AfZJ50ViC5
YZClYOLGv0zexWW71/Iht2ondEHIFv6nw5CvtIem9yglDIfF0BbRtGGzpRZH3Mfr/NvT2VfIu2IN
VeAN3t2YiWc9Je3OYkga18nnsqlrP1NL5cjdj0WHfx8Os8j5lwopSsaaKBeOSkO9DUrVcVhlepZs
mtM0aOWcY9E9xgJJuRlC1wfI13bfISXI7FoCrYPTZAhiudCEim4vcOL4tpj2NYqpGRaMDwx95ZEI
KuCs1f4q8X3vyVXb4PXfiSKTiOJYVtCgFICTjqJAz8RTBQWT+5Mz78luqcPSU5PEAJ6C4S+IFmie
Ariw2yk/MR8dFAOTqyBVBcaKOKmHH6b+JqpxwSiYIRZM+21pjmcKlXCIXRfFSHry1cPcUIXqBqK+
I9LPL6TUE25VlP0a9H+2iesd4+fg0E900A46jI2waIk1S6I6ihiJw2AGyLqzje/jt5vXsKseCZfk
rSDhQgNJj5ypFc8mhAqPTbgXtWn2xDVp9ZDWGL0GWuATdqZJJC4MOPfmwpIOQdShhkbj8xZ1w5lM
fPJTS4hrVpEZhqdZlZekXqiE98xc7qM3UQjUAIJfW9Ejj2vArmTp17q/0KdyRL4B2hsfqVV8SYHO
6/XE8Bm+pplylG+IBbsoa43yIDJ+y33VQfz5DUTXERitcSPcgJkSr2OhPWuwPhQQE6AQWbmSGhMQ
GIDQiVIljFWA3OyWZwS9oMWa2e9alVUEQG7f/LKbNZyzDbMKbgygriWwzi1tDqVae82Z0oJj8uDK
HmmoVZG/MO53WI3kTzPbvjO37hzVhQRTrQ/tsFQl3GLJn0Fts4sjgbO+aee8Pf22a9lMqzgxXMiM
ti9g73n66iVb3BTAiWx7s3o8xN36Xt4VBE2G49iwI0/hieHwdf2K5KrsBR7Y4rQGVT9w+6NukT2Q
Fia7zl8Km29KjIxrrvCAyUjZ7tak/u3NdFGbt/Dh0aj2gR9Yo4qAkeI0mNUOpLiQKpUt8BKIBWEj
5u0hN7cBuAmQIcmy/45jA6k8WBiEK3381b4VgG3ul0NhDj0LIE1BYuNn3iPedsylYcMCx14ZEPou
vGoGkrr5rIGi4MdSKXgpSTSMyxggZh/Cv5tLothMafaKq2bbpwDbDWyD+TwWe6/+FxK02s7MQgRy
ri0RbWhZp//sVLt9ZzxSV/8IMLJads+S8GPoB8HhIrJYa8tHe/p/RQLIlzQo0AelIQNH30rIjnNm
N7xszkgWVizNPWiSI7gM1QCFZrAfS7drkGvBBr2qdm6SJzeBPPyOweAHTs2cJ5FVo1MDXlzhWYf2
fjSNW+1lcAeOfvzpqX8V17KrqLvKC+FQ1Zf6K4rkheUa+TzHeVyWRaocdK+8goP1OFG1VR5I/j89
JHJhP0EAq1g2oH7DilYe945lMl4+dZhOFNUB1Zcd0scMpMyAHcp6cbaTuk6F1JULldfFmSA/BUQ/
oa66XpW/nNwTpb28Y5kgiGVo0UaUbFNSvWxzy+9zmDbiOymMMQTO6/XBuUVhY/U4DT7Styfqa34J
H39pSO5vLHqV7ObjlVwGlWqFo8ATl5PoCXY1WCxntWg2kCJThJQJw/lJVDxwubgqNNWRHNy/CcoS
1v+f6obIBYT3XYZCRa+MsDwODglW7bE2r0Vg0O5yVALr9cWtNt3Wk7QYyX/l9rjqgdfDFcSoyJ1P
hACMryrjvQfPxWSb1RLxpmKlFTj/EmiVCXyActwxI66desDP67HF7/l8nGYt/WL8VuwjlLCKOHnE
RaDf/CnXe8f11XuCmpJDgQTqiyC4gZ6o3CcvSM9IDmJAyP3z8uB2UUURg4vVSlVj1V1sYXj+ToTi
qzDiSrioJPlnJem7TVstThe0BQ4xrwaX0hkVFXyWWtAajhTN6JcsAN0extJo9vDdeO5hewq5ZJvr
1wf57EwpzgSaWf3rp5h8328jRCqBjoKdsOAi/tn6b90hxOuTvzi9C5qam7PWGjl7xaUT7Zj4ksyW
yw+/sX3HiJG7wYPhkq5vxGAEDMNEAacNGftzpiIIt4+oX0k5K4c9Iz9cTCWWfoYtJ4HZlf7nbC+A
cbEej0bV2ZEIAkIZ9DzE9MusDDSzs5sou3uflK8ZV3S4iWDb5qE1FW0+AP3uiimbVyAlCtG3aEGn
MtqM99w4vRZ0T0vdeg7nSVvDIf3FVH/VPg4VpgeSaCb1wJoi+F0jRMw39Xiq2YhCVnx7gwfxcy9P
b5YDQeCwjqWK/fTgmJO2kzi8QaSumm7p6QxWQWaN+kcNgHJJUq9QypopDaVXjyg+BVesD2ppq9NA
ylE03o26BWXS/9nsTQf6NZxvAa3MMsYWcs9OI+n0Mfl87fldYQ1YxbmZWoW+L+gJ6zIJFxFYDjNE
k1UtplgkENsXpVD7f/8P+7fy3tPUtb701x08Ow63afz0ty0u6yPZT963sn3TsJq/1u5bYg3jYj7S
jo6ayj1ePzqCb8KrDNPBXLCEj0Ryjl/e1v9Hu/k4/nEQWPNvX862bhGzINuLuZ0ggCn8ZvOGy+Rj
Nfe7eNmScfr6ZLW6vaJFsK/k9mu6sWZ2W2XRV3FPBrqv0RuKpgVFBAfd3XhSjjODddCij+ZWzOwM
MTzi37rSiQ5ivoQ/3XXOUJJlxVMH7igm4DziObN/YiNdKEd+j0WB4w1sFco8KEz7+dx5CGZXdZWB
3V0nIdUsMV4W8aCyF3fXeGOKVFTCwZ3aziLPsZoClMCnWY4uvvIedpUhr7Piz7rr2M9lEtwulPND
3tWku3JemdcYSU+85UQUpQ3rwbgv8xSWMeutXtiFYggUT+zEER4i/yEl6y53IgBMX3hXwSKXOJeF
1TMj7/HMeTzjFPnHVb7kvtZwKYTUKgho1b4OCwSyTJ2zh/JAK/U0FMgv9znBBtRGZMt2EPgHdfBC
2uCTwpL5ZDZyJRKcYPYQSRLYWCktfFKf09gOSG2tc3ZpeUhyUukXnJMaSlrMWZiZ0ADbE/bDe9Nn
3+Y1Q0mz2u4agMGA/O+BZoPHXPHAo9f2esdT/zSniMfyf+y2R2weqATDe+Ey7aECFy1src+5BVKx
9Q2ZZJz6KKcRHUQI83xMst4hsdUB9rK9go669oNeintVCFljpU65MO3loh5SJZzGzb6M7TXV5dVx
j386lpFVXCTTF/FRkWBb+aCnJ0EAqLsEaSttwYbhmR8vgQ4LFXXwIYuwelsLYCRWqs9zfsoWHVpu
987uct27rvZq3yAD1ddWFAIjgnXU2OANo1+SB1rqP7AbJ6rU9YHYuUgwG9xQ4yDkOHKIg+ZHWIRx
GgHTzvqTJMDSluHni3VxnPYz8O1/8G3FjGm71uljS/iEi6KLpGTEPOefSuJkBfiFjToK5uFCl44d
JBdytlymHbRmY53Zb9k690Swlw//KJoZ/dSM/EwPzM2KbJewkTg2+ArbrJh3eekodxRwKK5JvgtV
URGe5cNcKezu2cxGgICR0QYDL2WYVPBkVr+aCUba27kMujS9KLBJZMuMDVeZJVNwABwLre7P77yo
AU/1D+zU/O5r8g9mWLvr3za+Php/Y2Vw1hknfrBiWIoh1VupAiuaOi8WJinWji0SANbhmVpaaFJH
qX0EaTUAmdGtGhya2TYiDjKNyFAQyq8u2s64AzbkWYNduobS+Oezojmjyf1Y9vQIebU9grOi0rff
MXpJ3YvcZIAW56jUp4q8XX0QPfunLBNKAfeF5gudlxVzOdPxqESHGNGKDv6Pbue3ha4hCW9TbcPG
1Dy0L8hXcc+1LWgMt6swRmVUnWVInw1JI92bqFDwT9aik1GEd8YZPq6zCIGwQpvXUrRoIfAFshY4
URSxOru49be/eDFQv8f+27OsLl2xyLnuRqkdy0hdwRM3/pFzwpBKXBdLM9EnZ/VneT2JV1wGBD6P
PtKW05G7mXQ51F/amQkdTqSvEQVaDGjJTIhpATyVwemITTbRUFjdLhI0c9mHJ7AqDHz4ZOxD9BN/
y/1t+zpE7spvknR09EoLSZka4dQCCxWwaunRwFaaZPMMgq1HkyrUk7Xqp20/CIvC8TjwRXRD0gnq
1uaZBL9ysbEH65tcigxTlorrOTGal0q6SKEeKx6Kb/eA55AvINXD0+Qhs7kqSDn6v4e2vOgYrdvo
v7x03uf1xgy3BpJdEVY72kasjeB5ZnUVkTmAks1WRuXRJbgXf5JUpRlnrpE87qyc1p9EaA4RtFnh
6D4rpEb3+1HTtCFWTlUic2eJPiBYcA4dcA8j8LET+yfqU3a+MmhMHnZSvdFXsc/KEMK4yPJG4v5s
5dM+axaZDPyor2mswglkctNVTqCUTvltlSMaPOhlgjDl4pL2Y28/dK8XNx3TPmNXKQAU2BCfUPey
kmpX5mxqNSRzTpOmHYhugGc3k8bxRQRQ2G7Egydkoa/qoROQvuwlEd0J/8LfpsE53MK8skMRugtW
gHRF/03z/akVEk7bMKoH/4lFx6bqzZ1chSOnn0ql3NpQBn9VHlJtRHALskiRhsV8WL4vYP9d04US
fQi0DJdfkGjsr7GuY8tAEkIR6FKwAPHMBioTZcvyVPrsI5V9poCg4Vpb8JNLp1oxI5LPeSvGr2QQ
hr0UcH70O/gjDNKgYuslKUsv40XDHkvVbE9WopxGE0xhdCzON0PreLw7lSrrjZatj31ENGaYg/fp
kxhhJ9Gdrb9EDJhuXuvoGQuYjrBmVmR2woXQu5G45q2XhI9pL+HD/FjwGK+NGgnU1UwFNSlQW0vO
TZEdQMYxykpPRxI+IcibMDQ6o14Szg9d+2pNK/YpGru2xbissesCljS6V83kNTbExsowATNiW6yS
/z3k2y+d81rrQ3n/qmWtD9HuY/8Jh9DTzISxFLX6fm/3IrTNyUlSF3RvHrzpRtMtB7xav4rCu9AP
wvCS074WWpqtakcwnxuUCWjhrVL3BmbvxP+j+aWBGEUFshQSKlLPYAdho+bcQGXNnN7MhlPc43Kw
cLR/WoC6e+K6R6Fq1I3aysaQadWn5q5J5mgIWp3xQyuJefEGdM0JvJyQEx3HQn1fuEKYQDrpmDg6
X3mY6/cWNR8CHVnc4foSz9c7+lph0QS/W98uDaVgVS9KR0ssO6ouVoMetWz5HwawYJMn5C/jDzo8
eE5ib51Y1Se+JJhQsSLbqzmMWhzBobon8u1hgmifjS8QIqwOsOqU+b2lw/kApj71FMj1c3f8UxKl
qlJGrBxF55i+R6HvJ5jlDKXIakKGd3a1Ys+/Oe6OevHt1E/uD9jmU9vV1vOakwQmfxu+LxX0AtBF
7N3gIEHbidlD1fua75eOgnqW3VgZdtbFk+m+hpJH+bjXJhdcYY4xoZoeCjbnsavLZrtpCfIL5tgX
dkvPxZ6tKpzy2YmnOkcbvMY4hAYIPyZZRxGUaguO6XlJCm5UM08BtJtJOsMWvHI8c9Q0eNt37Pw5
8f/dhrGwDz31s/RzcuS/atlYUFUJ0+iYEYjyzpDTijQyLjoo3pq3gSNOZ2YSZVWEDvr60o2cvIX1
ThcsZk9Pom4KCg1Kt1yPG4EyHYCiQ+b1CCFM3KfeRMk5aiYFabq3t3PBSjGYMqlyBPMKlgF7tw91
WtHy1y502UiZRj8Kkzk+Ft1IA0Uqroq4S/Jgm9CPWZ7zOXZ2abScFVI2hNcDN7ZT5z6r44Nu/1eG
/hclAxJ9SIyYrDv19vCXrPvTJ4fU5UjUPGHr2fQBl6NeCnDW45TjgYOrcdRZ46eUcsyxGp7PVJ4a
Xcfx9LowvYr/K5oiImr/EYnMHQHZHTywKravdrYhGDbXSXTyHkBz3YHaLs8HEFcr0CxpK1NfGM6M
seKIpCtpJW0qnZ3an76M+0piY3s+l2FdP7OfmrvJyb3BkGkz4yE7Va6Vyg9k1+bbEcxljxeQglmX
fBZ6NJPsNEkLpf4JQMjQdGt1JfFGoryyC1MLureqAwcm3zS1aantHVvACgf7O+asYyYogS2ShyFr
0Pq9XcFGiTWnP+aYUeFdgpBXQmOk1RXnAkKZjgaC6H11SY7ReZ5Cdozp/WxgBZri8iLOaXTiRx/H
X7/W82FJWtO+3ePrTDEDgV9fT3qh3JWQYivInBY6p8m1avNVXWD5WZ4VXBPPXL8Q96T6D7Wp41cf
zICFyCtixgdtoACGJ0Pskp7fnIb7NQTorxFlnhh1HxsblwaDuSl/h8DyP7bcnz7Tf8y5LKSHfg8I
Zp/daoDIlJevrtcxcz42ggB6eEqSwG541WU+whTbk3rzCWKg/IhWESDWj5lDqCnpQiP8w5ETFiBk
sUFNFW4jGHeD6KJpDoMhbYYyeFd05xSmKzUlMsPGlDpatIklFmVtTc4hg7Ny9XhWiY+KzQEFOhc0
0LPRcPg8JdG7Xd/sbIBmIVNUUJTchwCzeM2fliVpgfRk1Lw6QQ1n6KcG3mUt6ZIfJur6gAlXN6SG
HDeiHxSaEbKU91RVCjqkJsBr6gRQDiZ1ZyayXXeCbcvOT5/SSDyAeQPfcL3Zeq2t1CWeYYhwjjng
sH9f+bGHzRaMA2aMjadpPoyfsx6I6sNgkJ6/7kVsHpvzURQozmSkq9v7NJvNkL3ZZNBrJjvHROLs
rUZQN/lI/v+Bf+ZIR5M5ylctjAWg3gj1kX+PWSUB6nA8nBFJLjUkt0Qy9cjaQkC4Dq932+hF0H5e
R1+BF8auJBYKAWAY3kUPTpVOg0t8mdroZ4yFHZN6ddyOoMjUus1nIxs8z3NZKQUDYrd3pTyzRfEM
9CUJR9OgFzHrwC/u+3NqydjvDE0yOaF6Advfmm/OnWvyBmOFYf1o9knVtZ115o5umgZEdb7giZ8x
jCbtk49J54IqmjGq7FVZ/kTKSgfWmIz/osTLC2dEfz/w76sWZwGvx9S8qVi8tgCTe2zXgZ4ANcMK
KjKdhE0ffH9p6pLYDLNp8H1Gdw8y3HHX0QTj2xAuN1ZJN403W4/N6OyJoo4H8589ncZXGgZYa+HV
+O8LiB93SnQtTCJS1GTvsCRZuTp2SwgBilviPDNNKyqhf3qNkgpYeMYVdT+d2Wvb8Hd5dZNHJ+4O
f8aLanJpEsFITrBA5KtDmFPfPv+aXvSY2RXkMYGEYwhpBQjl05YTxK6QrOHYQAYOtj/f9tLP6vYy
gldJny3uX5sM3yN1XUQgMTWST1vA/EO9y5QwncJRmhR4l0AjDp/F5qdHKb43aiCUDSx3NTmlM8bC
m3KOm+/bikuiC8W6JPIxA6jUsk27U8M=
`pragma protect end_protected
