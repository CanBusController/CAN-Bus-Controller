-- Network_can.vhd

-- Generated using ACDS version 13.1 162 at 2017.01.15.11:33:35

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity Network_can is
	port (
		clk_0_clk : in std_logic := '0'; -- clk_0.clk
		clk_clk   : in std_logic := '0'  --   clk.clk
	);
end entity Network_can;

architecture rtl of Network_can is
	component CAN_Controller_top is
		port (
			read      : in  std_logic                     := 'X';             -- read
			write     : in  std_logic                     := 'X';             -- write
			address   : in  std_logic_vector(5 downto 0)  := (others => 'X'); -- address
			writedata : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata  : out std_logic_vector(15 downto 0);                    -- readdata
			rst       : in  std_logic                     := 'X';             -- reset
			clk       : in  std_logic                     := 'X';             -- clk
			RxCAN     : in  std_logic                     := 'X';             -- export
			TxCAN     : out std_logic                                         -- export
		);
	end component CAN_Controller_top;

	component Network_can_nios2_qsys_0 is
		port (
			clk                                   : in  std_logic                     := 'X';             -- clk
			reset_n                               : in  std_logic                     := 'X';             -- reset_n
			reset_req                             : in  std_logic                     := 'X';             -- reset_req
			d_address                             : out std_logic_vector(13 downto 0);                    -- address
			d_byteenable                          : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                                : out std_logic;                                        -- read
			d_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			d_write                               : out std_logic;                                        -- write
			d_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_debug_module_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                             : out std_logic_vector(13 downto 0);                    -- address
			i_read                                : out std_logic;                                        -- read
			i_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			d_irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			jtag_debug_module_resetrequest        : out std_logic;                                        -- reset
			jtag_debug_module_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			jtag_debug_module_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			jtag_debug_module_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			jtag_debug_module_read                : in  std_logic                     := 'X';             -- read
			jtag_debug_module_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			jtag_debug_module_waitrequest         : out std_logic;                                        -- waitrequest
			jtag_debug_module_write               : in  std_logic                     := 'X';             -- write
			jtag_debug_module_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			no_ci_readra                          : out std_logic                                         -- readra
		);
	end component Network_can_nios2_qsys_0;

	component Network_can_nios2_qsys_1 is
		port (
			clk                                   : in  std_logic                     := 'X';             -- clk
			reset_n                               : in  std_logic                     := 'X';             -- reset_n
			reset_req                             : in  std_logic                     := 'X';             -- reset_req
			d_address                             : out std_logic_vector(13 downto 0);                    -- address
			d_byteenable                          : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                                : out std_logic;                                        -- read
			d_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			d_write                               : out std_logic;                                        -- write
			d_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_debug_module_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                             : out std_logic_vector(13 downto 0);                    -- address
			i_read                                : out std_logic;                                        -- read
			i_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			d_irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			jtag_debug_module_resetrequest        : out std_logic;                                        -- reset
			jtag_debug_module_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			jtag_debug_module_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			jtag_debug_module_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			jtag_debug_module_read                : in  std_logic                     := 'X';             -- read
			jtag_debug_module_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			jtag_debug_module_waitrequest         : out std_logic;                                        -- waitrequest
			jtag_debug_module_write               : in  std_logic                     := 'X';             -- write
			jtag_debug_module_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			no_ci_readra                          : out std_logic                                         -- readra
		);
	end component Network_can_nios2_qsys_1;

	component Network_can_onchip_memory2_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(10 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X'              -- reset_req
		);
	end component Network_can_onchip_memory2_0;

	component Network_can_onchip_memory2_1 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(10 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X'              -- reset_req
		);
	end component Network_can_onchip_memory2_1;

	component can_BUS is
		port (
			rx1 : out std_logic;        -- export
			tx1 : in  std_logic := 'X'; -- export
			rx2 : out std_logic;        -- export
			tx2 : in  std_logic := 'X'  -- export
		);
	end component can_BUS;

	component Network_can_mm_interconnect_0 is
		port (
			clk_0_clk_clk                                    : in  std_logic                     := 'X';             -- clk
			nios2_qsys_0_reset_n_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			nios2_qsys_0_data_master_address                 : in  std_logic_vector(13 downto 0) := (others => 'X'); -- address
			nios2_qsys_0_data_master_waitrequest             : out std_logic;                                        -- waitrequest
			nios2_qsys_0_data_master_byteenable              : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			nios2_qsys_0_data_master_read                    : in  std_logic                     := 'X';             -- read
			nios2_qsys_0_data_master_readdata                : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_qsys_0_data_master_write                   : in  std_logic                     := 'X';             -- write
			nios2_qsys_0_data_master_writedata               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			nios2_qsys_0_data_master_debugaccess             : in  std_logic                     := 'X';             -- debugaccess
			nios2_qsys_0_instruction_master_address          : in  std_logic_vector(13 downto 0) := (others => 'X'); -- address
			nios2_qsys_0_instruction_master_waitrequest      : out std_logic;                                        -- waitrequest
			nios2_qsys_0_instruction_master_read             : in  std_logic                     := 'X';             -- read
			nios2_qsys_0_instruction_master_readdata         : out std_logic_vector(31 downto 0);                    -- readdata
			Can_controller_0_avalon_slave_0_address          : out std_logic_vector(5 downto 0);                     -- address
			Can_controller_0_avalon_slave_0_write            : out std_logic;                                        -- write
			Can_controller_0_avalon_slave_0_read             : out std_logic;                                        -- read
			Can_controller_0_avalon_slave_0_readdata         : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			Can_controller_0_avalon_slave_0_writedata        : out std_logic_vector(15 downto 0);                    -- writedata
			nios2_qsys_0_jtag_debug_module_address           : out std_logic_vector(8 downto 0);                     -- address
			nios2_qsys_0_jtag_debug_module_write             : out std_logic;                                        -- write
			nios2_qsys_0_jtag_debug_module_read              : out std_logic;                                        -- read
			nios2_qsys_0_jtag_debug_module_readdata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios2_qsys_0_jtag_debug_module_writedata         : out std_logic_vector(31 downto 0);                    -- writedata
			nios2_qsys_0_jtag_debug_module_byteenable        : out std_logic_vector(3 downto 0);                     -- byteenable
			nios2_qsys_0_jtag_debug_module_waitrequest       : in  std_logic                     := 'X';             -- waitrequest
			nios2_qsys_0_jtag_debug_module_debugaccess       : out std_logic;                                        -- debugaccess
			onchip_memory2_0_s1_address                      : out std_logic_vector(10 downto 0);                    -- address
			onchip_memory2_0_s1_write                        : out std_logic;                                        -- write
			onchip_memory2_0_s1_readdata                     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			onchip_memory2_0_s1_writedata                    : out std_logic_vector(15 downto 0);                    -- writedata
			onchip_memory2_0_s1_byteenable                   : out std_logic_vector(1 downto 0);                     -- byteenable
			onchip_memory2_0_s1_chipselect                   : out std_logic;                                        -- chipselect
			onchip_memory2_0_s1_clken                        : out std_logic                                         -- clken
		);
	end component Network_can_mm_interconnect_0;

	component Network_can_mm_interconnect_1 is
		port (
			clk_1_clk_clk                                    : in  std_logic                     := 'X';             -- clk
			nios2_qsys_1_reset_n_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			nios2_qsys_1_data_master_address                 : in  std_logic_vector(13 downto 0) := (others => 'X'); -- address
			nios2_qsys_1_data_master_waitrequest             : out std_logic;                                        -- waitrequest
			nios2_qsys_1_data_master_byteenable              : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			nios2_qsys_1_data_master_read                    : in  std_logic                     := 'X';             -- read
			nios2_qsys_1_data_master_readdata                : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_qsys_1_data_master_write                   : in  std_logic                     := 'X';             -- write
			nios2_qsys_1_data_master_writedata               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			nios2_qsys_1_data_master_debugaccess             : in  std_logic                     := 'X';             -- debugaccess
			nios2_qsys_1_instruction_master_address          : in  std_logic_vector(13 downto 0) := (others => 'X'); -- address
			nios2_qsys_1_instruction_master_waitrequest      : out std_logic;                                        -- waitrequest
			nios2_qsys_1_instruction_master_read             : in  std_logic                     := 'X';             -- read
			nios2_qsys_1_instruction_master_readdata         : out std_logic_vector(31 downto 0);                    -- readdata
			Can_controller_1_avalon_slave_0_address          : out std_logic_vector(5 downto 0);                     -- address
			Can_controller_1_avalon_slave_0_write            : out std_logic;                                        -- write
			Can_controller_1_avalon_slave_0_read             : out std_logic;                                        -- read
			Can_controller_1_avalon_slave_0_readdata         : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			Can_controller_1_avalon_slave_0_writedata        : out std_logic_vector(15 downto 0);                    -- writedata
			nios2_qsys_1_jtag_debug_module_address           : out std_logic_vector(8 downto 0);                     -- address
			nios2_qsys_1_jtag_debug_module_write             : out std_logic;                                        -- write
			nios2_qsys_1_jtag_debug_module_read              : out std_logic;                                        -- read
			nios2_qsys_1_jtag_debug_module_readdata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios2_qsys_1_jtag_debug_module_writedata         : out std_logic_vector(31 downto 0);                    -- writedata
			nios2_qsys_1_jtag_debug_module_byteenable        : out std_logic_vector(3 downto 0);                     -- byteenable
			nios2_qsys_1_jtag_debug_module_waitrequest       : in  std_logic                     := 'X';             -- waitrequest
			nios2_qsys_1_jtag_debug_module_debugaccess       : out std_logic;                                        -- debugaccess
			onchip_memory2_1_s1_address                      : out std_logic_vector(10 downto 0);                    -- address
			onchip_memory2_1_s1_write                        : out std_logic;                                        -- write
			onchip_memory2_1_s1_readdata                     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			onchip_memory2_1_s1_writedata                    : out std_logic_vector(15 downto 0);                    -- writedata
			onchip_memory2_1_s1_byteenable                   : out std_logic_vector(1 downto 0);                     -- byteenable
			onchip_memory2_1_s1_chipselect                   : out std_logic;                                        -- chipselect
			onchip_memory2_1_s1_clken                        : out std_logic                                         -- clken
		);
	end component Network_can_mm_interconnect_1;

	component Network_can_irq_mapper is
		port (
			clk        : in  std_logic                     := 'X'; -- clk
			reset      : in  std_logic                     := 'X'; -- reset
			sender_irq : out std_logic_vector(31 downto 0)         -- irq
		);
	end component Network_can_irq_mapper;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			reset_in1      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal nios2_qsys_0_jtag_debug_module_reset_reset                   : std_logic;                     -- nios2_qsys_0:jtag_debug_module_resetrequest -> [rst_controller:reset_in0, rst_controller:reset_in1]
	signal nios2_qsys_1_jtag_debug_module_reset_reset                   : std_logic;                     -- nios2_qsys_1:jtag_debug_module_resetrequest -> [rst_controller_001:reset_in0, rst_controller_001:reset_in1]
	signal bus_can_0_conduit_end_export                                 : std_logic;                     -- Bus_CAN_0:rx1 -> Can_controller_0:RxCAN
	signal can_controller_0_conduit_end_1_export                        : std_logic;                     -- Can_controller_0:TxCAN -> Bus_CAN_0:tx1
	signal bus_can_0_conduit_end_2_export                               : std_logic;                     -- Bus_CAN_0:rx2 -> Can_controller_1:RxCAN
	signal can_controller_1_conduit_end_1_export                        : std_logic;                     -- Can_controller_1:TxCAN -> Bus_CAN_0:tx2
	signal nios2_qsys_0_data_master_waitrequest                         : std_logic;                     -- mm_interconnect_0:nios2_qsys_0_data_master_waitrequest -> nios2_qsys_0:d_waitrequest
	signal nios2_qsys_0_data_master_writedata                           : std_logic_vector(31 downto 0); -- nios2_qsys_0:d_writedata -> mm_interconnect_0:nios2_qsys_0_data_master_writedata
	signal nios2_qsys_0_data_master_address                             : std_logic_vector(13 downto 0); -- nios2_qsys_0:d_address -> mm_interconnect_0:nios2_qsys_0_data_master_address
	signal nios2_qsys_0_data_master_write                               : std_logic;                     -- nios2_qsys_0:d_write -> mm_interconnect_0:nios2_qsys_0_data_master_write
	signal nios2_qsys_0_data_master_read                                : std_logic;                     -- nios2_qsys_0:d_read -> mm_interconnect_0:nios2_qsys_0_data_master_read
	signal nios2_qsys_0_data_master_readdata                            : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_qsys_0_data_master_readdata -> nios2_qsys_0:d_readdata
	signal nios2_qsys_0_data_master_debugaccess                         : std_logic;                     -- nios2_qsys_0:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:nios2_qsys_0_data_master_debugaccess
	signal nios2_qsys_0_data_master_byteenable                          : std_logic_vector(3 downto 0);  -- nios2_qsys_0:d_byteenable -> mm_interconnect_0:nios2_qsys_0_data_master_byteenable
	signal mm_interconnect_0_onchip_memory2_0_s1_writedata              : std_logic_vector(15 downto 0); -- mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	signal mm_interconnect_0_onchip_memory2_0_s1_address                : std_logic_vector(10 downto 0); -- mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	signal mm_interconnect_0_onchip_memory2_0_s1_chipselect             : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	signal mm_interconnect_0_onchip_memory2_0_s1_clken                  : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	signal mm_interconnect_0_onchip_memory2_0_s1_write                  : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	signal mm_interconnect_0_onchip_memory2_0_s1_readdata               : std_logic_vector(15 downto 0); -- onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	signal mm_interconnect_0_onchip_memory2_0_s1_byteenable             : std_logic_vector(1 downto 0);  -- mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	signal nios2_qsys_0_instruction_master_waitrequest                  : std_logic;                     -- mm_interconnect_0:nios2_qsys_0_instruction_master_waitrequest -> nios2_qsys_0:i_waitrequest
	signal nios2_qsys_0_instruction_master_address                      : std_logic_vector(13 downto 0); -- nios2_qsys_0:i_address -> mm_interconnect_0:nios2_qsys_0_instruction_master_address
	signal nios2_qsys_0_instruction_master_read                         : std_logic;                     -- nios2_qsys_0:i_read -> mm_interconnect_0:nios2_qsys_0_instruction_master_read
	signal nios2_qsys_0_instruction_master_readdata                     : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_qsys_0_instruction_master_readdata -> nios2_qsys_0:i_readdata
	signal mm_interconnect_0_can_controller_0_avalon_slave_0_writedata  : std_logic_vector(15 downto 0); -- mm_interconnect_0:Can_controller_0_avalon_slave_0_writedata -> Can_controller_0:writedata
	signal mm_interconnect_0_can_controller_0_avalon_slave_0_address    : std_logic_vector(5 downto 0);  -- mm_interconnect_0:Can_controller_0_avalon_slave_0_address -> Can_controller_0:address
	signal mm_interconnect_0_can_controller_0_avalon_slave_0_write      : std_logic;                     -- mm_interconnect_0:Can_controller_0_avalon_slave_0_write -> Can_controller_0:write
	signal mm_interconnect_0_can_controller_0_avalon_slave_0_read       : std_logic;                     -- mm_interconnect_0:Can_controller_0_avalon_slave_0_read -> Can_controller_0:read
	signal mm_interconnect_0_can_controller_0_avalon_slave_0_readdata   : std_logic_vector(15 downto 0); -- Can_controller_0:readdata -> mm_interconnect_0:Can_controller_0_avalon_slave_0_readdata
	signal mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest : std_logic;                     -- nios2_qsys_0:jtag_debug_module_waitrequest -> mm_interconnect_0:nios2_qsys_0_jtag_debug_module_waitrequest
	signal mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata   : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_qsys_0_jtag_debug_module_writedata -> nios2_qsys_0:jtag_debug_module_writedata
	signal mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address     : std_logic_vector(8 downto 0);  -- mm_interconnect_0:nios2_qsys_0_jtag_debug_module_address -> nios2_qsys_0:jtag_debug_module_address
	signal mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write       : std_logic;                     -- mm_interconnect_0:nios2_qsys_0_jtag_debug_module_write -> nios2_qsys_0:jtag_debug_module_write
	signal mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read        : std_logic;                     -- mm_interconnect_0:nios2_qsys_0_jtag_debug_module_read -> nios2_qsys_0:jtag_debug_module_read
	signal mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata    : std_logic_vector(31 downto 0); -- nios2_qsys_0:jtag_debug_module_readdata -> mm_interconnect_0:nios2_qsys_0_jtag_debug_module_readdata
	signal mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess : std_logic;                     -- mm_interconnect_0:nios2_qsys_0_jtag_debug_module_debugaccess -> nios2_qsys_0:jtag_debug_module_debugaccess
	signal mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable  : std_logic_vector(3 downto 0);  -- mm_interconnect_0:nios2_qsys_0_jtag_debug_module_byteenable -> nios2_qsys_0:jtag_debug_module_byteenable
	signal mm_interconnect_1_nios2_qsys_1_jtag_debug_module_waitrequest : std_logic;                     -- nios2_qsys_1:jtag_debug_module_waitrequest -> mm_interconnect_1:nios2_qsys_1_jtag_debug_module_waitrequest
	signal mm_interconnect_1_nios2_qsys_1_jtag_debug_module_writedata   : std_logic_vector(31 downto 0); -- mm_interconnect_1:nios2_qsys_1_jtag_debug_module_writedata -> nios2_qsys_1:jtag_debug_module_writedata
	signal mm_interconnect_1_nios2_qsys_1_jtag_debug_module_address     : std_logic_vector(8 downto 0);  -- mm_interconnect_1:nios2_qsys_1_jtag_debug_module_address -> nios2_qsys_1:jtag_debug_module_address
	signal mm_interconnect_1_nios2_qsys_1_jtag_debug_module_write       : std_logic;                     -- mm_interconnect_1:nios2_qsys_1_jtag_debug_module_write -> nios2_qsys_1:jtag_debug_module_write
	signal mm_interconnect_1_nios2_qsys_1_jtag_debug_module_read        : std_logic;                     -- mm_interconnect_1:nios2_qsys_1_jtag_debug_module_read -> nios2_qsys_1:jtag_debug_module_read
	signal mm_interconnect_1_nios2_qsys_1_jtag_debug_module_readdata    : std_logic_vector(31 downto 0); -- nios2_qsys_1:jtag_debug_module_readdata -> mm_interconnect_1:nios2_qsys_1_jtag_debug_module_readdata
	signal mm_interconnect_1_nios2_qsys_1_jtag_debug_module_debugaccess : std_logic;                     -- mm_interconnect_1:nios2_qsys_1_jtag_debug_module_debugaccess -> nios2_qsys_1:jtag_debug_module_debugaccess
	signal mm_interconnect_1_nios2_qsys_1_jtag_debug_module_byteenable  : std_logic_vector(3 downto 0);  -- mm_interconnect_1:nios2_qsys_1_jtag_debug_module_byteenable -> nios2_qsys_1:jtag_debug_module_byteenable
	signal mm_interconnect_1_can_controller_1_avalon_slave_0_writedata  : std_logic_vector(15 downto 0); -- mm_interconnect_1:Can_controller_1_avalon_slave_0_writedata -> Can_controller_1:writedata
	signal mm_interconnect_1_can_controller_1_avalon_slave_0_address    : std_logic_vector(5 downto 0);  -- mm_interconnect_1:Can_controller_1_avalon_slave_0_address -> Can_controller_1:address
	signal mm_interconnect_1_can_controller_1_avalon_slave_0_write      : std_logic;                     -- mm_interconnect_1:Can_controller_1_avalon_slave_0_write -> Can_controller_1:write
	signal mm_interconnect_1_can_controller_1_avalon_slave_0_read       : std_logic;                     -- mm_interconnect_1:Can_controller_1_avalon_slave_0_read -> Can_controller_1:read
	signal mm_interconnect_1_can_controller_1_avalon_slave_0_readdata   : std_logic_vector(15 downto 0); -- Can_controller_1:readdata -> mm_interconnect_1:Can_controller_1_avalon_slave_0_readdata
	signal nios2_qsys_1_instruction_master_waitrequest                  : std_logic;                     -- mm_interconnect_1:nios2_qsys_1_instruction_master_waitrequest -> nios2_qsys_1:i_waitrequest
	signal nios2_qsys_1_instruction_master_address                      : std_logic_vector(13 downto 0); -- nios2_qsys_1:i_address -> mm_interconnect_1:nios2_qsys_1_instruction_master_address
	signal nios2_qsys_1_instruction_master_read                         : std_logic;                     -- nios2_qsys_1:i_read -> mm_interconnect_1:nios2_qsys_1_instruction_master_read
	signal nios2_qsys_1_instruction_master_readdata                     : std_logic_vector(31 downto 0); -- mm_interconnect_1:nios2_qsys_1_instruction_master_readdata -> nios2_qsys_1:i_readdata
	signal mm_interconnect_1_onchip_memory2_1_s1_writedata              : std_logic_vector(15 downto 0); -- mm_interconnect_1:onchip_memory2_1_s1_writedata -> onchip_memory2_1:writedata
	signal mm_interconnect_1_onchip_memory2_1_s1_address                : std_logic_vector(10 downto 0); -- mm_interconnect_1:onchip_memory2_1_s1_address -> onchip_memory2_1:address
	signal mm_interconnect_1_onchip_memory2_1_s1_chipselect             : std_logic;                     -- mm_interconnect_1:onchip_memory2_1_s1_chipselect -> onchip_memory2_1:chipselect
	signal mm_interconnect_1_onchip_memory2_1_s1_clken                  : std_logic;                     -- mm_interconnect_1:onchip_memory2_1_s1_clken -> onchip_memory2_1:clken
	signal mm_interconnect_1_onchip_memory2_1_s1_write                  : std_logic;                     -- mm_interconnect_1:onchip_memory2_1_s1_write -> onchip_memory2_1:write
	signal mm_interconnect_1_onchip_memory2_1_s1_readdata               : std_logic_vector(15 downto 0); -- onchip_memory2_1:readdata -> mm_interconnect_1:onchip_memory2_1_s1_readdata
	signal mm_interconnect_1_onchip_memory2_1_s1_byteenable             : std_logic_vector(1 downto 0);  -- mm_interconnect_1:onchip_memory2_1_s1_byteenable -> onchip_memory2_1:byteenable
	signal nios2_qsys_1_data_master_waitrequest                         : std_logic;                     -- mm_interconnect_1:nios2_qsys_1_data_master_waitrequest -> nios2_qsys_1:d_waitrequest
	signal nios2_qsys_1_data_master_writedata                           : std_logic_vector(31 downto 0); -- nios2_qsys_1:d_writedata -> mm_interconnect_1:nios2_qsys_1_data_master_writedata
	signal nios2_qsys_1_data_master_address                             : std_logic_vector(13 downto 0); -- nios2_qsys_1:d_address -> mm_interconnect_1:nios2_qsys_1_data_master_address
	signal nios2_qsys_1_data_master_write                               : std_logic;                     -- nios2_qsys_1:d_write -> mm_interconnect_1:nios2_qsys_1_data_master_write
	signal nios2_qsys_1_data_master_read                                : std_logic;                     -- nios2_qsys_1:d_read -> mm_interconnect_1:nios2_qsys_1_data_master_read
	signal nios2_qsys_1_data_master_readdata                            : std_logic_vector(31 downto 0); -- mm_interconnect_1:nios2_qsys_1_data_master_readdata -> nios2_qsys_1:d_readdata
	signal nios2_qsys_1_data_master_debugaccess                         : std_logic;                     -- nios2_qsys_1:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_1:nios2_qsys_1_data_master_debugaccess
	signal nios2_qsys_1_data_master_byteenable                          : std_logic_vector(3 downto 0);  -- nios2_qsys_1:d_byteenable -> mm_interconnect_1:nios2_qsys_1_data_master_byteenable
	signal nios2_qsys_0_d_irq_irq                                       : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> nios2_qsys_0:d_irq
	signal nios2_qsys_1_d_irq_irq                                       : std_logic_vector(31 downto 0); -- irq_mapper_001:sender_irq -> nios2_qsys_1:d_irq
	signal rst_controller_reset_out_reset                               : std_logic;                     -- rst_controller:reset_out -> [Can_controller_0:rst, irq_mapper:reset, mm_interconnect_0:nios2_qsys_0_reset_n_reset_bridge_in_reset_reset, onchip_memory2_0:reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                           : std_logic;                     -- rst_controller:reset_req -> [nios2_qsys_0:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	signal rst_controller_001_reset_out_reset                           : std_logic;                     -- rst_controller_001:reset_out -> [Can_controller_1:rst, irq_mapper_001:reset, mm_interconnect_1:nios2_qsys_1_reset_n_reset_bridge_in_reset_reset, onchip_memory2_1:reset, rst_controller_001_reset_out_reset:in, rst_translator_001:in_reset]
	signal rst_controller_001_reset_out_reset_req                       : std_logic;                     -- rst_controller_001:reset_req -> [nios2_qsys_1:reset_req, onchip_memory2_1:reset_req, rst_translator_001:reset_req_in]
	signal rst_controller_reset_out_reset_ports_inv                     : std_logic;                     -- rst_controller_reset_out_reset:inv -> nios2_qsys_0:reset_n
	signal rst_controller_001_reset_out_reset_ports_inv                 : std_logic;                     -- rst_controller_001_reset_out_reset:inv -> nios2_qsys_1:reset_n

begin

	can_controller_0 : component CAN_Controller_top
		port map (
			read      => mm_interconnect_0_can_controller_0_avalon_slave_0_read,      -- avalon_slave_0.read
			write     => mm_interconnect_0_can_controller_0_avalon_slave_0_write,     --               .write
			address   => mm_interconnect_0_can_controller_0_avalon_slave_0_address,   --               .address
			writedata => mm_interconnect_0_can_controller_0_avalon_slave_0_writedata, --               .writedata
			readdata  => mm_interconnect_0_can_controller_0_avalon_slave_0_readdata,  --               .readdata
			rst       => rst_controller_reset_out_reset,                              --     reset_sink.reset
			clk       => clk_clk,                                                     --     clock_sink.clk
			RxCAN     => bus_can_0_conduit_end_export,                                --    conduit_end.export
			TxCAN     => can_controller_0_conduit_end_1_export                        --  conduit_end_1.export
		);

	nios2_qsys_0 : component Network_can_nios2_qsys_0
		port map (
			clk                                   => clk_clk,                                                      --                       clk.clk
			reset_n                               => rst_controller_reset_out_reset_ports_inv,                     --                   reset_n.reset_n
			reset_req                             => rst_controller_reset_out_reset_req,                           --                          .reset_req
			d_address                             => nios2_qsys_0_data_master_address,                             --               data_master.address
			d_byteenable                          => nios2_qsys_0_data_master_byteenable,                          --                          .byteenable
			d_read                                => nios2_qsys_0_data_master_read,                                --                          .read
			d_readdata                            => nios2_qsys_0_data_master_readdata,                            --                          .readdata
			d_waitrequest                         => nios2_qsys_0_data_master_waitrequest,                         --                          .waitrequest
			d_write                               => nios2_qsys_0_data_master_write,                               --                          .write
			d_writedata                           => nios2_qsys_0_data_master_writedata,                           --                          .writedata
			jtag_debug_module_debugaccess_to_roms => nios2_qsys_0_data_master_debugaccess,                         --                          .debugaccess
			i_address                             => nios2_qsys_0_instruction_master_address,                      --        instruction_master.address
			i_read                                => nios2_qsys_0_instruction_master_read,                         --                          .read
			i_readdata                            => nios2_qsys_0_instruction_master_readdata,                     --                          .readdata
			i_waitrequest                         => nios2_qsys_0_instruction_master_waitrequest,                  --                          .waitrequest
			d_irq                                 => nios2_qsys_0_d_irq_irq,                                       --                     d_irq.irq
			jtag_debug_module_resetrequest        => nios2_qsys_0_jtag_debug_module_reset_reset,                   --   jtag_debug_module_reset.reset
			jtag_debug_module_address             => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address,     --         jtag_debug_module.address
			jtag_debug_module_byteenable          => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable,  --                          .byteenable
			jtag_debug_module_debugaccess         => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess, --                          .debugaccess
			jtag_debug_module_read                => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read,        --                          .read
			jtag_debug_module_readdata            => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata,    --                          .readdata
			jtag_debug_module_waitrequest         => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest, --                          .waitrequest
			jtag_debug_module_write               => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write,       --                          .write
			jtag_debug_module_writedata           => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata,   --                          .writedata
			no_ci_readra                          => open                                                          -- custom_instruction_master.readra
		);

	nios2_qsys_1 : component Network_can_nios2_qsys_1
		port map (
			clk                                   => clk_0_clk,                                                    --                       clk.clk
			reset_n                               => rst_controller_001_reset_out_reset_ports_inv,                 --                   reset_n.reset_n
			reset_req                             => rst_controller_001_reset_out_reset_req,                       --                          .reset_req
			d_address                             => nios2_qsys_1_data_master_address,                             --               data_master.address
			d_byteenable                          => nios2_qsys_1_data_master_byteenable,                          --                          .byteenable
			d_read                                => nios2_qsys_1_data_master_read,                                --                          .read
			d_readdata                            => nios2_qsys_1_data_master_readdata,                            --                          .readdata
			d_waitrequest                         => nios2_qsys_1_data_master_waitrequest,                         --                          .waitrequest
			d_write                               => nios2_qsys_1_data_master_write,                               --                          .write
			d_writedata                           => nios2_qsys_1_data_master_writedata,                           --                          .writedata
			jtag_debug_module_debugaccess_to_roms => nios2_qsys_1_data_master_debugaccess,                         --                          .debugaccess
			i_address                             => nios2_qsys_1_instruction_master_address,                      --        instruction_master.address
			i_read                                => nios2_qsys_1_instruction_master_read,                         --                          .read
			i_readdata                            => nios2_qsys_1_instruction_master_readdata,                     --                          .readdata
			i_waitrequest                         => nios2_qsys_1_instruction_master_waitrequest,                  --                          .waitrequest
			d_irq                                 => nios2_qsys_1_d_irq_irq,                                       --                     d_irq.irq
			jtag_debug_module_resetrequest        => nios2_qsys_1_jtag_debug_module_reset_reset,                   --   jtag_debug_module_reset.reset
			jtag_debug_module_address             => mm_interconnect_1_nios2_qsys_1_jtag_debug_module_address,     --         jtag_debug_module.address
			jtag_debug_module_byteenable          => mm_interconnect_1_nios2_qsys_1_jtag_debug_module_byteenable,  --                          .byteenable
			jtag_debug_module_debugaccess         => mm_interconnect_1_nios2_qsys_1_jtag_debug_module_debugaccess, --                          .debugaccess
			jtag_debug_module_read                => mm_interconnect_1_nios2_qsys_1_jtag_debug_module_read,        --                          .read
			jtag_debug_module_readdata            => mm_interconnect_1_nios2_qsys_1_jtag_debug_module_readdata,    --                          .readdata
			jtag_debug_module_waitrequest         => mm_interconnect_1_nios2_qsys_1_jtag_debug_module_waitrequest, --                          .waitrequest
			jtag_debug_module_write               => mm_interconnect_1_nios2_qsys_1_jtag_debug_module_write,       --                          .write
			jtag_debug_module_writedata           => mm_interconnect_1_nios2_qsys_1_jtag_debug_module_writedata,   --                          .writedata
			no_ci_readra                          => open                                                          -- custom_instruction_master.readra
		);

	onchip_memory2_0 : component Network_can_onchip_memory2_0
		port map (
			clk        => clk_clk,                                          --   clk1.clk
			address    => mm_interconnect_0_onchip_memory2_0_s1_address,    --     s1.address
			clken      => mm_interconnect_0_onchip_memory2_0_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_onchip_memory2_0_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_onchip_memory2_0_s1_write,      --       .write
			readdata   => mm_interconnect_0_onchip_memory2_0_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_onchip_memory2_0_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_onchip_memory2_0_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,                   -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req                --       .reset_req
		);

	onchip_memory2_1 : component Network_can_onchip_memory2_1
		port map (
			clk        => clk_0_clk,                                        --   clk1.clk
			address    => mm_interconnect_1_onchip_memory2_1_s1_address,    --     s1.address
			clken      => mm_interconnect_1_onchip_memory2_1_s1_clken,      --       .clken
			chipselect => mm_interconnect_1_onchip_memory2_1_s1_chipselect, --       .chipselect
			write      => mm_interconnect_1_onchip_memory2_1_s1_write,      --       .write
			readdata   => mm_interconnect_1_onchip_memory2_1_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_1_onchip_memory2_1_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_1_onchip_memory2_1_s1_byteenable, --       .byteenable
			reset      => rst_controller_001_reset_out_reset,               -- reset1.reset
			reset_req  => rst_controller_001_reset_out_reset_req            --       .reset_req
		);

	can_controller_1 : component CAN_Controller_top
		port map (
			read      => mm_interconnect_1_can_controller_1_avalon_slave_0_read,      -- avalon_slave_0.read
			write     => mm_interconnect_1_can_controller_1_avalon_slave_0_write,     --               .write
			address   => mm_interconnect_1_can_controller_1_avalon_slave_0_address,   --               .address
			writedata => mm_interconnect_1_can_controller_1_avalon_slave_0_writedata, --               .writedata
			readdata  => mm_interconnect_1_can_controller_1_avalon_slave_0_readdata,  --               .readdata
			rst       => rst_controller_001_reset_out_reset,                          --     reset_sink.reset
			clk       => clk_0_clk,                                                   --     clock_sink.clk
			RxCAN     => bus_can_0_conduit_end_2_export,                              --    conduit_end.export
			TxCAN     => can_controller_1_conduit_end_1_export                        --  conduit_end_1.export
		);

	bus_can_0 : component can_BUS
		port map (
			rx1 => bus_can_0_conduit_end_export,          --   conduit_end.export
			tx1 => can_controller_0_conduit_end_1_export, -- conduit_end_1.export
			rx2 => bus_can_0_conduit_end_2_export,        -- conduit_end_2.export
			tx2 => can_controller_1_conduit_end_1_export  -- conduit_end_3.export
		);

	mm_interconnect_0 : component Network_can_mm_interconnect_0
		port map (
			clk_0_clk_clk                                    => clk_clk,                                                      --                                  clk_0_clk.clk
			nios2_qsys_0_reset_n_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                               -- nios2_qsys_0_reset_n_reset_bridge_in_reset.reset
			nios2_qsys_0_data_master_address                 => nios2_qsys_0_data_master_address,                             --                   nios2_qsys_0_data_master.address
			nios2_qsys_0_data_master_waitrequest             => nios2_qsys_0_data_master_waitrequest,                         --                                           .waitrequest
			nios2_qsys_0_data_master_byteenable              => nios2_qsys_0_data_master_byteenable,                          --                                           .byteenable
			nios2_qsys_0_data_master_read                    => nios2_qsys_0_data_master_read,                                --                                           .read
			nios2_qsys_0_data_master_readdata                => nios2_qsys_0_data_master_readdata,                            --                                           .readdata
			nios2_qsys_0_data_master_write                   => nios2_qsys_0_data_master_write,                               --                                           .write
			nios2_qsys_0_data_master_writedata               => nios2_qsys_0_data_master_writedata,                           --                                           .writedata
			nios2_qsys_0_data_master_debugaccess             => nios2_qsys_0_data_master_debugaccess,                         --                                           .debugaccess
			nios2_qsys_0_instruction_master_address          => nios2_qsys_0_instruction_master_address,                      --            nios2_qsys_0_instruction_master.address
			nios2_qsys_0_instruction_master_waitrequest      => nios2_qsys_0_instruction_master_waitrequest,                  --                                           .waitrequest
			nios2_qsys_0_instruction_master_read             => nios2_qsys_0_instruction_master_read,                         --                                           .read
			nios2_qsys_0_instruction_master_readdata         => nios2_qsys_0_instruction_master_readdata,                     --                                           .readdata
			Can_controller_0_avalon_slave_0_address          => mm_interconnect_0_can_controller_0_avalon_slave_0_address,    --            Can_controller_0_avalon_slave_0.address
			Can_controller_0_avalon_slave_0_write            => mm_interconnect_0_can_controller_0_avalon_slave_0_write,      --                                           .write
			Can_controller_0_avalon_slave_0_read             => mm_interconnect_0_can_controller_0_avalon_slave_0_read,       --                                           .read
			Can_controller_0_avalon_slave_0_readdata         => mm_interconnect_0_can_controller_0_avalon_slave_0_readdata,   --                                           .readdata
			Can_controller_0_avalon_slave_0_writedata        => mm_interconnect_0_can_controller_0_avalon_slave_0_writedata,  --                                           .writedata
			nios2_qsys_0_jtag_debug_module_address           => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address,     --             nios2_qsys_0_jtag_debug_module.address
			nios2_qsys_0_jtag_debug_module_write             => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write,       --                                           .write
			nios2_qsys_0_jtag_debug_module_read              => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read,        --                                           .read
			nios2_qsys_0_jtag_debug_module_readdata          => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata,    --                                           .readdata
			nios2_qsys_0_jtag_debug_module_writedata         => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata,   --                                           .writedata
			nios2_qsys_0_jtag_debug_module_byteenable        => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable,  --                                           .byteenable
			nios2_qsys_0_jtag_debug_module_waitrequest       => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest, --                                           .waitrequest
			nios2_qsys_0_jtag_debug_module_debugaccess       => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess, --                                           .debugaccess
			onchip_memory2_0_s1_address                      => mm_interconnect_0_onchip_memory2_0_s1_address,                --                        onchip_memory2_0_s1.address
			onchip_memory2_0_s1_write                        => mm_interconnect_0_onchip_memory2_0_s1_write,                  --                                           .write
			onchip_memory2_0_s1_readdata                     => mm_interconnect_0_onchip_memory2_0_s1_readdata,               --                                           .readdata
			onchip_memory2_0_s1_writedata                    => mm_interconnect_0_onchip_memory2_0_s1_writedata,              --                                           .writedata
			onchip_memory2_0_s1_byteenable                   => mm_interconnect_0_onchip_memory2_0_s1_byteenable,             --                                           .byteenable
			onchip_memory2_0_s1_chipselect                   => mm_interconnect_0_onchip_memory2_0_s1_chipselect,             --                                           .chipselect
			onchip_memory2_0_s1_clken                        => mm_interconnect_0_onchip_memory2_0_s1_clken                   --                                           .clken
		);

	mm_interconnect_1 : component Network_can_mm_interconnect_1
		port map (
			clk_1_clk_clk                                    => clk_0_clk,                                                    --                                  clk_1_clk.clk
			nios2_qsys_1_reset_n_reset_bridge_in_reset_reset => rst_controller_001_reset_out_reset,                           -- nios2_qsys_1_reset_n_reset_bridge_in_reset.reset
			nios2_qsys_1_data_master_address                 => nios2_qsys_1_data_master_address,                             --                   nios2_qsys_1_data_master.address
			nios2_qsys_1_data_master_waitrequest             => nios2_qsys_1_data_master_waitrequest,                         --                                           .waitrequest
			nios2_qsys_1_data_master_byteenable              => nios2_qsys_1_data_master_byteenable,                          --                                           .byteenable
			nios2_qsys_1_data_master_read                    => nios2_qsys_1_data_master_read,                                --                                           .read
			nios2_qsys_1_data_master_readdata                => nios2_qsys_1_data_master_readdata,                            --                                           .readdata
			nios2_qsys_1_data_master_write                   => nios2_qsys_1_data_master_write,                               --                                           .write
			nios2_qsys_1_data_master_writedata               => nios2_qsys_1_data_master_writedata,                           --                                           .writedata
			nios2_qsys_1_data_master_debugaccess             => nios2_qsys_1_data_master_debugaccess,                         --                                           .debugaccess
			nios2_qsys_1_instruction_master_address          => nios2_qsys_1_instruction_master_address,                      --            nios2_qsys_1_instruction_master.address
			nios2_qsys_1_instruction_master_waitrequest      => nios2_qsys_1_instruction_master_waitrequest,                  --                                           .waitrequest
			nios2_qsys_1_instruction_master_read             => nios2_qsys_1_instruction_master_read,                         --                                           .read
			nios2_qsys_1_instruction_master_readdata         => nios2_qsys_1_instruction_master_readdata,                     --                                           .readdata
			Can_controller_1_avalon_slave_0_address          => mm_interconnect_1_can_controller_1_avalon_slave_0_address,    --            Can_controller_1_avalon_slave_0.address
			Can_controller_1_avalon_slave_0_write            => mm_interconnect_1_can_controller_1_avalon_slave_0_write,      --                                           .write
			Can_controller_1_avalon_slave_0_read             => mm_interconnect_1_can_controller_1_avalon_slave_0_read,       --                                           .read
			Can_controller_1_avalon_slave_0_readdata         => mm_interconnect_1_can_controller_1_avalon_slave_0_readdata,   --                                           .readdata
			Can_controller_1_avalon_slave_0_writedata        => mm_interconnect_1_can_controller_1_avalon_slave_0_writedata,  --                                           .writedata
			nios2_qsys_1_jtag_debug_module_address           => mm_interconnect_1_nios2_qsys_1_jtag_debug_module_address,     --             nios2_qsys_1_jtag_debug_module.address
			nios2_qsys_1_jtag_debug_module_write             => mm_interconnect_1_nios2_qsys_1_jtag_debug_module_write,       --                                           .write
			nios2_qsys_1_jtag_debug_module_read              => mm_interconnect_1_nios2_qsys_1_jtag_debug_module_read,        --                                           .read
			nios2_qsys_1_jtag_debug_module_readdata          => mm_interconnect_1_nios2_qsys_1_jtag_debug_module_readdata,    --                                           .readdata
			nios2_qsys_1_jtag_debug_module_writedata         => mm_interconnect_1_nios2_qsys_1_jtag_debug_module_writedata,   --                                           .writedata
			nios2_qsys_1_jtag_debug_module_byteenable        => mm_interconnect_1_nios2_qsys_1_jtag_debug_module_byteenable,  --                                           .byteenable
			nios2_qsys_1_jtag_debug_module_waitrequest       => mm_interconnect_1_nios2_qsys_1_jtag_debug_module_waitrequest, --                                           .waitrequest
			nios2_qsys_1_jtag_debug_module_debugaccess       => mm_interconnect_1_nios2_qsys_1_jtag_debug_module_debugaccess, --                                           .debugaccess
			onchip_memory2_1_s1_address                      => mm_interconnect_1_onchip_memory2_1_s1_address,                --                        onchip_memory2_1_s1.address
			onchip_memory2_1_s1_write                        => mm_interconnect_1_onchip_memory2_1_s1_write,                  --                                           .write
			onchip_memory2_1_s1_readdata                     => mm_interconnect_1_onchip_memory2_1_s1_readdata,               --                                           .readdata
			onchip_memory2_1_s1_writedata                    => mm_interconnect_1_onchip_memory2_1_s1_writedata,              --                                           .writedata
			onchip_memory2_1_s1_byteenable                   => mm_interconnect_1_onchip_memory2_1_s1_byteenable,             --                                           .byteenable
			onchip_memory2_1_s1_chipselect                   => mm_interconnect_1_onchip_memory2_1_s1_chipselect,             --                                           .chipselect
			onchip_memory2_1_s1_clken                        => mm_interconnect_1_onchip_memory2_1_s1_clken                   --                                           .clken
		);

	irq_mapper : component Network_can_irq_mapper
		port map (
			clk        => clk_clk,                        --       clk.clk
			reset      => rst_controller_reset_out_reset, -- clk_reset.reset
			sender_irq => nios2_qsys_0_d_irq_irq          --    sender.irq
		);

	irq_mapper_001 : component Network_can_irq_mapper
		port map (
			clk        => clk_0_clk,                          --       clk.clk
			reset      => rst_controller_001_reset_out_reset, -- clk_reset.reset
			sender_irq => nios2_qsys_1_d_irq_irq              --    sender.irq
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => nios2_qsys_0_jtag_debug_module_reset_reset, -- reset_in0.reset
			reset_in1      => nios2_qsys_0_jtag_debug_module_reset_reset, -- reset_in1.reset
			clk            => clk_clk,                                    --       clk.clk
			reset_out      => rst_controller_reset_out_reset,             -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req,         --          .reset_req
			reset_req_in0  => '0',                                        -- (terminated)
			reset_req_in1  => '0',                                        -- (terminated)
			reset_in2      => '0',                                        -- (terminated)
			reset_req_in2  => '0',                                        -- (terminated)
			reset_in3      => '0',                                        -- (terminated)
			reset_req_in3  => '0',                                        -- (terminated)
			reset_in4      => '0',                                        -- (terminated)
			reset_req_in4  => '0',                                        -- (terminated)
			reset_in5      => '0',                                        -- (terminated)
			reset_req_in5  => '0',                                        -- (terminated)
			reset_in6      => '0',                                        -- (terminated)
			reset_req_in6  => '0',                                        -- (terminated)
			reset_in7      => '0',                                        -- (terminated)
			reset_req_in7  => '0',                                        -- (terminated)
			reset_in8      => '0',                                        -- (terminated)
			reset_req_in8  => '0',                                        -- (terminated)
			reset_in9      => '0',                                        -- (terminated)
			reset_req_in9  => '0',                                        -- (terminated)
			reset_in10     => '0',                                        -- (terminated)
			reset_req_in10 => '0',                                        -- (terminated)
			reset_in11     => '0',                                        -- (terminated)
			reset_req_in11 => '0',                                        -- (terminated)
			reset_in12     => '0',                                        -- (terminated)
			reset_req_in12 => '0',                                        -- (terminated)
			reset_in13     => '0',                                        -- (terminated)
			reset_req_in13 => '0',                                        -- (terminated)
			reset_in14     => '0',                                        -- (terminated)
			reset_req_in14 => '0',                                        -- (terminated)
			reset_in15     => '0',                                        -- (terminated)
			reset_req_in15 => '0'                                         -- (terminated)
		);

	rst_controller_001 : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => nios2_qsys_1_jtag_debug_module_reset_reset, -- reset_in0.reset
			reset_in1      => nios2_qsys_1_jtag_debug_module_reset_reset, -- reset_in1.reset
			clk            => clk_0_clk,                                  --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset,         -- reset_out.reset
			reset_req      => rst_controller_001_reset_out_reset_req,     --          .reset_req
			reset_req_in0  => '0',                                        -- (terminated)
			reset_req_in1  => '0',                                        -- (terminated)
			reset_in2      => '0',                                        -- (terminated)
			reset_req_in2  => '0',                                        -- (terminated)
			reset_in3      => '0',                                        -- (terminated)
			reset_req_in3  => '0',                                        -- (terminated)
			reset_in4      => '0',                                        -- (terminated)
			reset_req_in4  => '0',                                        -- (terminated)
			reset_in5      => '0',                                        -- (terminated)
			reset_req_in5  => '0',                                        -- (terminated)
			reset_in6      => '0',                                        -- (terminated)
			reset_req_in6  => '0',                                        -- (terminated)
			reset_in7      => '0',                                        -- (terminated)
			reset_req_in7  => '0',                                        -- (terminated)
			reset_in8      => '0',                                        -- (terminated)
			reset_req_in8  => '0',                                        -- (terminated)
			reset_in9      => '0',                                        -- (terminated)
			reset_req_in9  => '0',                                        -- (terminated)
			reset_in10     => '0',                                        -- (terminated)
			reset_req_in10 => '0',                                        -- (terminated)
			reset_in11     => '0',                                        -- (terminated)
			reset_req_in11 => '0',                                        -- (terminated)
			reset_in12     => '0',                                        -- (terminated)
			reset_req_in12 => '0',                                        -- (terminated)
			reset_in13     => '0',                                        -- (terminated)
			reset_req_in13 => '0',                                        -- (terminated)
			reset_in14     => '0',                                        -- (terminated)
			reset_req_in14 => '0',                                        -- (terminated)
			reset_in15     => '0',                                        -- (terminated)
			reset_req_in15 => '0'                                         -- (terminated)
		);

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

end architecture rtl; -- of Network_can
