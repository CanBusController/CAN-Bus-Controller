// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
eAUqrAONsFa09d64yFz192HN2oYdp7/NvgTSdQtDo98CbVtgQa6Z38DT/GQHg2WUQOVDkTVbBLyR
vAZzSQgYwh1VYnFT4N6QLssda1XkpcEgmoB6dqMwA9QH4C+bwW/zzou7NDlOwNX132ISsrtZOeHl
Oae5vAj28mYJUJxjGzTt0hiCXpOH4nKtxbRtzqNsPiXPvN0cyqZsJpbrVcQrl5QHATjXBK+tTpMB
04ozmcR2aABBP2Yh3p239WnADDJcT8UB8BIS7KoDjjzNcdAX8yDQFuKSvCij3vzXVcaCruWxDUTf
wkN7jkS2jYX6Z/yGl1EoWNIOQb9U3y7Nbjka2w==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
4aD5XzEsdl97f4VMDB/h9GVmQskrvdMlEytegrcC0sXVuk4FG7wJKtXYQdVYeKXBOoIljrs454VH
GnUoFjj46I15XIMRZw9c4TpqoQGOn/7oukaD3XLTU6M8Rb6f0PCA2KtbnmVySsxm45O/Q9Id0qOO
Ae7x0P8cawlTvLCx8LjpvnssZJjBvflJmM3/Hk/3nrKOTV+GHsYPV2Hmxfj7ntEE8nCCWf4aLMbl
reqfRGU0/IarUO25ldOlQQB7uUCgw9MzMVS4psx+zRH2RLL/z6gfrs3sQiMWMkOHjfyol0nKLhni
8GuRJQ3/Vl2wOAMGEcx1aLaRRBhuIwZwrcZmj7iciPgO9aN/rK7wJkv2fYMDoYNU1oR9HL3rTcnk
nz9V4rMJw+weEAB1t4UWRyBSevfzyc560wuASMh3a9d8SYNux99bpAPG2v75YJWwp4by0wUzXD/D
I7AN1aZrTKku8hLfPYUNr+AkGJyaSDE49dobK7DOM1sURJLbQqdXzKMNHahbzpqGpv9/G9ipsgiJ
F3PIS8Vz884Bn5rKAJ6S9GZfACXSCwXJJBm3y6ip0ZCAkGExKpucaedowQfOlLCHYVKxkw2AVLOb
qX9C+4l28m5rExOLT6pmEa7RxPDJ0ZyZKkuv4oXhVDD9c66tuqRR83itA5s5cNqOtYMDcqXl4oo4
+58m2RYlEXViAwAvpnUVysiWuNv5jqMsd2RUTrdyTv05xRSV1se/MmW3t8PV7ngl8+aIXHGZsAjJ
68/OUYF6BmZoxBD55f7TLu8O48IHnIgbOFjOLuhBYqXtaYdmWxM7uZy2zm5+J8sw8z0qxpEkAWK4
ntIAaKkP2vqyABhEm9nANr/ba9K4/bB52oh0VcVCR36Ti1H1UcnHki04eKrIpneSiksRNvHipd+n
uJ4Z/hfZ2JUSIRjswbNWY8BPQoIw8pr57f2NmdzWanAUBASwAJrz57QBjJbnMCf61YvOnly0MDP/
e7g/hMZfvTyGNmMAZ0yzv5XVncFokA9iEsrCQZaan5+MXho/nN2xlbP2H/Ehhh4PS0eqnDsX8Gjm
sIqIFGfBmT5zHASYoiLC+eumYUfTZ4ktAhu9V06sCpL8SV7lHserCm6E0WoDnqy5S2wGeOubYvHC
6AYNMa5m1Jl1ZsxVoJW2e9hZb/nFxTQCpkDbjsDzCJQ72LehG4mZrWeVXLHNqO7NFpDn4ZOP3tKZ
RjH2kjwIJITfiEQP3CDa0SCF8sFqQe/NuTbV2lLSmPZQiHF+ST79dWxHw5G/JSNKRJQH/FfUBSEI
gnw0SqGYY4PRC5yW/Bq35YKWyUR7D8uB4XVMl6OkTK1ljgUfllMUfWylPApZpJIWO4FTEyIjsjJ5
uZ16iQNdDymPll4JDioqyzlHMsiEGkGSrggeAteGxMzkv6kgp7ZwIUgEXXXyyzCd96UCIVnN5Nts
9MUcsu8NmnfF0wDQYcGRfpPX8KRs7hok56Ou1x9YaX+Asf7d/jIxkxt4io9trNRcDwoEbXNcBrLf
WgEbzKzciUMVtZMESmcuY0OKOt+a0TE1L6P9EiArx1TfWNKFaWWsRgAPabXk98HWaUttZ1JAWHIi
Gs0QYxZOJLmUuHvd5ElgXzECYuIDpBv+st8X8JrUtNnmj0VzukKMic0dy9otE5+eNTJ0bxo0l36m
XleVlarUOEOWP77exAAlruC0jzLY7uqgYFoAaGIxnbwrVLWZf5JIHDT04jyJkNJTET1TaLTLFVBb
Piixk05F840p49r6jTYpgtuFjkE4Yvs1r/HuvNvJc8Tz/HqtqDrp7/NelUtIePvfHd1yaebBJzAm
uP/ZIoxWKtiSZR7KoBUAeK3tCSMoqZePexk87ZHsHyxW7Dpjtbiuujz+2BhNqA4PzNuQ/Wr/98ql
poNeO/PmaxjxKQhj8BLcXRG0bS7YYSsPiGKCNArGZ4XSc25q8pQw9OGqy4sYb3VatSU/2PY7Rvfu
nbc+H1A+I3bN7bnHS59LgXmaZKRfa6NFx2Z2csab8q2hhibouRN+i5gF8a0nPBpLHqHo3YZXyb6N
1TavoY6wsh0YZuIRvetkGtNPiJT8UcI944HprDW+PWTHmia+zXsONIzvMrFyjHVd77Ho1eTeGydX
ld23hgJz6og4DNpHfYNaHtzRW1WktGaUIJRkX9MBKKQYBKSKx+ukB9vKr7rroy5UXe8ZPjXPf5GU
b/vpaQtmFKLnQ1JT/IBM1wJCRQxfmxdEtPba5N6ufknbf6a+Z1lmN29SUHGZzv2pQLPG42XvsaX2
ZEknyFigp/Wu17gV2d4y96P/up7TwAL0rvW2gU2rIVbZc9ga+P0nQ0M+eTcmJbe+9oJnHo74sxy/
/nBdX6mkJHjbu+6uJ/10SS53j6iI4PBTDeJzBJAb6+vF9/hrJKJdLR8XFN5Ub3ZTht7YFjdJBtVv
2J4g5VvpPXUwFovuvMGNnyG5Q89RJ+5jmeRWLiMPMl+kvw6T+2sfv551pcV4kboIDZxHZvH7h436
AZXgI5vJmvi6s78ASuo+5LF+M1r0WuY2eLQ3nflGhJpcM0AvdC7/P6dTwhb536YqgPi+006W3YgE
xq7YHQiqrGFmo7I7K9ff5z0u0lpyS/Qh4lVT+QsHGVV2BxdXCGoiSkejLZKtVntVQf0ybXd4hEb2
k06/f3z6hKJpITz9nhxTDlz6PvDhy6XrhpOKL3AzyMNZQoBO/AiJ6u6EF9tokzr063Z7Eij5kWjU
VCH34NnEH5bwvEhzM3CI5YBb3mszUoIG6DYF4mfsXLq0mlN4cfhGtX7CUGz6/A8LYE2WzshRGleL
Y6okkUbKt1VO3HtvUB4CXUvZZUX68kDhKZ0tZHTFYdnQtv+ata8mNQ0HRMZTMsTs4O7jcOUbzkw/
BRbmep2Itrhxza4lGYrsZKyDbioYmZljaEudKVPrdSm1P10aS+iopSFOgwzLOV7irTCVHbmcHSH2
oNSrP0R7ydsfq18mTl65CnJKHyfDBKMqTBuGNQn1rUwxSfzWFpD+X4S5yxtGEbMWRjFDCin9APRv
a9Mk4XzNzg8A4Zg7mwgc3uSy12PteE8Tx/ItCknMZxBZRwn9P2TkQ58AcsgCt2jty2Kcm0AXY5Ui
i6+2qOtnqSl4kh1g1jreQ0aJ+aTokXONyzjvIjqvdCGRG5o4I29JqSHb5l4RtM+XvgdihjOv4nsF
ZbPiakkZ+JybwZlh+ZtPft4dl1XPqDAdgSCBprMeWP8EkVQ+gXZl1zYzRFcY7/+HrTc7k5kf7COj
GoseDVXrDrEVhLi2I2ZdKzkVkA3Un0qX7+oArswWLIzRcjr+tf1ARs96/vBf2kN9ENy/S7C21/Hd
pkpmu7COgIltE2MsIBxqOIg43cK6j/lC6VJtYXn45Qcui5cMSSfGtk7vfhaBNb7bzXC8m4VyVjZ9
O55XbGgdp1DpXy+BlmQ21QpHZp5D+ly3YAOghnuCh4vccKwd+e04nzjOBqSgpRAz+/zTiqtObuES
zTMVR39PL2eOqnVIyMrbZruM01nYQFO3Ml9E00fZsi2gjLXJSZawDZtVDgGX6cPWwzR+QA1IYreM
j0HFPygxxA+Yi1OXQmqfoLYIBPCte+yIi7h0TKuQJDz3f9vXWLrM26HaZCrXdo+7U7bk6XlBweiD
k3JAXkn6vFary3eD97iGZ402fFkl9+avKefHO1/tEZTs752iSTFBsLMS3Z0a2wbKOeAJMHH3NR9J
FFGTb61EceBqIZng24qOBz0beCk4UNKgLVQwOgKy6zkQN2bU3KHucwqtoTA6d30HOPl/CTTseYtc
0AqdDRk40z3v1Wip0kMgSmB160uMKdMNdqGg8annCzyPPSuVdkczzg4tmJHW194nhV9ZZjGtxAgf
VactDUTWaJtc1Sth8M2r0lXa52/4onFnfUoQPLRFxH1kCSMZNxRzdmb7SjFv6yHe/eo+oB01zU/q
3FWczCIJ4v6rwTWSTnVePHofdeKJVmM3t0ffzz7R/2+ovfr/sPfSs3sRkTNKg4jda9puLolziedL
fBRToH6gmKX9u6OXslIMi5ZeTb4tZfbp4dKZvcQohd9RljnwGAR/YlTOoByqFO0me6ZHPnFg9qfz
hr9ZO6CJ+p1aZydwtAEdQX0fXY52MwyvVH0eCt72hrmAHjKvpU5lMR94aCKY1zzDPi94hKam4BkX
RrERjDG9vmDnZVYdEQgpYZYE3aI95i5W4RCO15ajJgef7I6pUdjy5GyAxw0IZIt8Fd5kvTFxUgKJ
oz02DFnUVCdyarDw+zinASk0rX/ChBCOrCIfArJ0DdqUoO+PEFfsz4oV/Y+z98bk5qbqk/kY5UxT
FBte/8DIEJLsSZLBWhICjfAY1qrq2ILFkq4ph88m+AkfHC4fPUPtOYwRlBef4fR9pPSP72beNRlk
F4ZRIdz5QS4NqrazURO6HcaKrXu4AuehFz+jmF+QmPM+rnbdZ8G/ZNsjbqxFHakOd/JM51JSPlnX
Px0Y2+/Jl+T6zxwjL6w9xhd3tQRy1JzR1VcJOfeNJ2GDZmjLIE6nWhobtOXeIrC1B4/DA9hT8VN+
as2eI0eeOOvFprR+bwI35xcaygaYU14fBKFAfc3ubUbVmwoEv9Dl4QRQDxqhDGXIeVoYOug1GtaA
1pReSZG3ApW6Bskbvb+A8ZmhV6UAY2Y7B3HB1soqTCjLwGXeDxbpONTh8NhVh3v9KuAN2GG+Mike
O8a1UiKxePh1I9MPDPjVRqhzFh9P7M8LlkVN1v+x+KBCY9OlBdrHlzAdGzN9+gj7tB8rYD19lk4t
wVuPjHIIHrc38zf3m+T+eg3u6+kbilPTIjo8rJXaxaxTHNx8seg3a3DvVueloAZy/NbbZXZW6J1+
SRqIYiDPxxZ0e9SzNu/ycSKKZ+oaJgZ70cyaFmu/holgEdjH3PPImJssLn8Ae/gnIha7EqL8rvqD
Cu7xYi+I5WgoKUI6tS1TuphfrRww2/ofu3a43t5713L2qaBExRvbHg6gWlLKiBINVKBHQULNODSP
K9hfqBaNqmUu3qPXfxRdPUsCgNzlaRblqeov4rgq08fLTvxjIxU8o4/UkFaXFxFLTyVF6TI47Cyl
PpbJ52dRZu8g4r2Pq+wzRXPSbTx1tFEXfRalMASwjjbZd8nvyjyEydlq5axmWLex9gYvAbhfK5bf
HvOWZe+3lo4yMxvy6b+EKPw45UpXYP5sBPVuwqFe1QcfXpLn7DgXkNTcy+OddKuh5bhhpKrV4huJ
NqFXKc3pdbw2DVnZYOUAFwRXcRRch/bqeZAmW7Td6M8ZiU3bWNaCVXuCtgQjvZqAfWXrhRFOTaup
pMdrPosqYUamhIX77pEqCk/0alfNOd8iyhNlLgNMevGf/OMMXLqqwWLN7MHERLsuq67uzv9pxa3A
ULCSUYmUkVvbdsBCF+sJ8Kh0hzRF9b9s8gTMF9TmzIoPVGP1bbnLpwqWkbUBlePXheQV2eaBICed
FZQ140R4RkqEnB1uFpzumWXxSgPXX1g3sTL2+HjYoKkf4bQUFJJ+dJXPu9RLZLXqZue3By0DfaCY
SpBCtbAGks3a0qnbgWXP/CFa12pkEYa77X83HtKmEKLJ3DZ/cUd7jzjNEaeZPmtRBQwj29ST6ePy
KWOIL0q7aFWqmltVjnMLpY5tQiuQzy3daBk7xiOGJoabKH+/uAf2RCu7+KoFn8itgUP/FifH3l5q
zSskKwoQRRgWKP5Ztq3MLCm9RBrCDg65XOKXOc/e2gz9y9J3+svL7xFgXfKaQqY9sAL0mxbIc6bu
Prd0+wSoRsT3EDrlx19GGgUbh5ByspuKCJNvXRkKWYpLtRpsUR0RAG10OLljiVDREEqWCCy0ZykB
QqsQjQZYDVZwBijCVBUhvm42+pEFxzpSrVYZEtCXZPfpV1pfF96s0qqiJp14ZUU7FYXNTotAg9EB
XJcoSF84JwTX/oXmjqKYL2AlTiSRSX169wa9MZPPW0QmXZVjR1g3xiw2nx9nvuwyuLuWDfCzqBer
9LvJrzJypjHIvRUMh9CrPTiyQkzhbU/04P3JNm9Cm28RpZky3b8kJyS7Xn9Y2rbV6jccEtcPYc2y
UEl4lmgP7BtaTpMBRitc5u3QbcucUapl/KGE01L3nU60yruD5l9OfHGGfQVEVpzBcF9qn0XJG8vT
L9NXnk0xYht1GZTetoUU9sPfV3mkrRIP6iPzS+Kjwv2lsLs0C1c/MtjtXBIeiHXF0CiZ7i10Fpt9
gMwJHVy8CsNOCMqBGZshYEgR7XnXGqOiWZum6lOQfnNSqGUY0ND7u/YPgKOOb/dSKOQWuIuw98HJ
RxEAjJiVqN162wbZHxY5k0xf//KhxOil2uIO4JsPVW8ZHrpZRX0Tq86VFMTnDvAeO+amyLtY6f6F
c8PYICRe9BDO9JTp3P8Dq8Oe7TsVtSV3COndVpVkrxjA9kgHzQBvYXOS1FqzeJba39VTtY0SnLrT
6Zyjj0HVVKDJQaPrlToWKqgxiuUmcc2vApxfyzlCqoviGI8Ig3WfMMUT0Zd4TlaMC/cbwqr0dQrG
MI4qlRJg9tynek+aK2irvDXZmTjUYrzZTzKvaJQ2Lsd0fFdDX23FaUy/7dw1nLTz0eL/e4Hzyj7M
TjXKQkTxjmRiwsTJ5Lj64DuptWv7ohVykB6mj1ITMiMTXa2saRMglw27v4nHJjD+mBP7/hVy86T3
ruCNeQ/Dd1mspnGcxgZNASbAwu4VgAbxXOnD4tacjwD+SmQNS55p21WRTSZnZyisNtxVAZ1anPkt
oV8kkZYj6x7/7kYc0q9EhuO+T7uMxljGHRJYOp4J/qFubCr6gkh0YmXrCHZxchScrxP+TD6/7ZfQ
kSGO29LWX5EVHRCaEkZR0HuvgEBwO/9ruuh93e0bs2yssY3w1kWUFbe1JGdGpOw7FL0DweDRgN0p
+xb8QjqIw5uq46mfqkwWkKQnbMgykqun56IFjwrYOybT7XWveDrrcmdWfNYZnbFlvculjvC6LoRt
LfNQNIMPtF/r3Nd7LyYye8CsMYWm2txcEVryY6psJxhscB5P8IUyMM4Pe7aIdQxQqQ6nAlfhJKFJ
V8FMT7PQfVDJDtyp5UQp9X7q+OzNPdIaGASRdP7OACeQBUY6om/aWKNUVusYoVvGxG8kuOxg3qZM
FcwacwKTdmyMPVU5ueyx/b/Bceurg2jiL/SzLDZ7vIxUUoX/WIHgy0NqqyghFMhoIlXBd+IpFxNK
1CEhdH3kurkT/AUHNzOcyh/2KnmUoQJqpry4fTlNXrVmJdRkOmwgDLhVDAP1V9FGI9m9RBi7mLaH
uVZgw0+4AhsVKhdIWvBQOiwQexFy95wrsr4IGpIrthJQDRqDG/F9Vb9DstHcX6mnlTGeuiqx80Vg
h+W9TZT9uE5eL2RO3Nmy2+yqGtflE5XHRAFrx42UGDECDq3WBKzfbQh8ambtoNESFQxoBq/NwIz8
L5lCoOi7qRa/2uOD2eNuqOYTcx2OvXTK1XoAby1Vt7h0+WfVNqKNWe89rQRZ24fhAFl4t6hvspa9
kFwDSU3Ru+bNsilEDa9mlpgC0rtzcdTgVLy/I5XbkYocQcUu16fGOuwFOicEd0V6A/sZM1ppwQji
if1vylKJryEZdlH2TXTAUWIBWyJj5HCNKl7cFZeDOOOKcY2pO4HSBL02HNHbat1Jqi6JWqlfyd5b
E+LW0M4N78oIODjv6L8pX/f+VgQiZIbujzja5hYHkvwD+HeSWX8/l3huS7PYuhCqKidGs5XbApYN
FB7nl8FawW0esINJkPcydVS8QtJ9XPPw3wr9XGFmoQJSuOUh+ps1s6JeCf9O5a/AYINSx+fHPEVa
j3pibULj1Tav3odJkT/tL2Tl99fuAtsNZRnTzbSQRRM7mqLfVxDmVwbNuDI/MbwM6Wm3HGndDZKw
7yHnGBWt5zkUcg78ODcDL4y0wBh0PQxU5DWiUjZkv+x7MhmAZ/7xKx4EG5fyidybIn9tpqpQR1ir
uqUCzHxrg1Gx7/42BesVeDfXgog+jmHtwz2D7Ksq/uk36ll+xI9CYdI/E/p7EhJgJXcD+Oo68YOB
boHKacbA2jcYkJbUUEZ4kXrKi8rf2Rl3QWk2yeYU53I7ygV/lD7/3cF5f10dBlfnAtFzzx4m09FY
8mWyVk/t3G80QahE/pGjVS4IRVBdLZw3+Za+/8U6Xl5e7KJX6l/Dybpqpxuq0qnzC/Sr+Se37bde
y6PrdNKwVj0N+JZoJUTwZx2pUmkHQh6MgYb9JigaoZ1UrLkpHYWmcczfOGqzE2rE8543WljR0aRj
NcRbYKo5/69U2Bw8oR7Ec9995mtpUbDTiQxiuJdUQtLjWi+t+24234+IxDBYXq+KGWuqJbIysYxI
VYrSEM65nuOQa6B77dl2Hw6DgL9oKNbqplO1wPpANAuA8PEL8eUr8EZ+ygP4JsvFjg6H0Xp4ZahI
erDbvSZQdigHUBMWSXL193+QQFzFMOHWQNbdYHSMZ657sLil6ykbdD5624cTRuylA/eZSGMRCobF
pkg/x+1WsKRw6yJntiT/x4BVz3kNQOiicinOqzFdhMpxorDcc8X8optwpQwQ7EwoC3DMGNhkg4ro
NQd/zuDXIZ8A4WTSW6yBTrZzfFKb4eWCyhSOsoqkBW+ENIeCy09EP5e/6g7Y7/jyUrKJ1bMvzmlT
pQs7P+Ji4qDUsDBVa48YvBXD5JxzRsbVo5zMA/27s8dQw0ajWnK7CCWe449U31d/qHEGz9fwFcfW
g4Wh+tTF/kwzqmptTx+2eXcNdrID21a0yp7eYK1Sg+hl6c17dWaXBzncg1H/V/0WnXqSZ35U70hq
x3huqBNdQHDbdZ010Cr7A0F/se6ye/DJbUerE3iPZoAnE8oHx+7+wKuZXkFSbkZ6MdvO6Bg1boZy
2bKTTPO+l7h3dhC7SGGFqIYozu7COn22fS5FJscIZXeJrNWd3VS6Ru2ftM1OFm7UXDXiF9l+8nAq
brSQol8NMUM5WDZEXXqY0bM5LHZIu5EFVzcaCpbH+6rbnJXTOwoT6h0hODq0KmLqO+c2CqES6Xae
0WHZSAejmvX1Un25MmesNSkRDpoSVm+zf9j3vP0U//mcPx2RNjsONJ4psYcV1bA4J0XLlSXIowQ0
EK+sQS6n2EfVg5w1PBa3HYA/vLqYeYOOWVh9z2s7SW/htvCgJiadQmF5MQ8wXq4RcC5wbh1pIkTU
PTRHAWJt+daEIBpXXLb6EctMFJGGI2TVaJSBbmP1K0z+Z0uJCQSbCK6PYrVy7hjjJJNpbQkVq+zy
wJC9mfKIqbqXyYZICISOPLTwF3bKWkgi6RAOt/teOY5SRTyGKW4cQ7XA1fS1OJpUvEUMRU8cwGm2
s6mEOE+vR8JnreSjCnp/K3xhr5klk38mSAn6wORUU0+kIMw+NDRkxtld1fP7USWFffgsC8UJcYlQ
Qu56ObdK2zFFqx21LcEbwcgdofAOxNESqJog4K2bbcoeBtRXfl+NBMJ+TTRT5XViaRNgg5nyuVju
tFcg/3hj5auPCdQou0AL0dk9W3sCOMl110kgdpsIwevJGKjQtKEHTRNDbcQELh6nDEvkwZMu0teU
l7bmvPcXBVFoqW4JR81PwI4LAJBujcKha00/ggl3hc0+sld/L9l2jnhsVAlmKwSUGMDcEzp+DI8P
5qeDOowDZV2cABAKabP4V8ojPaXr+hJggXhLzlwEfZUtwLYmovHqw+eYbE+OyVN1U37QiygrsGky
iX0yF/b5q/wfTnkx0s4o7jjOnqLtNAny3guwJJN07S7tiaFhtBsR+0EnLMm6mkS+nbV5H6WKpHF6
XMGcpMKdSqPFYvG+n5UFUnGn416jVPCHiHzrV8NkUI4kVf5r+bh5LDS4YdHElm9Oq11YIiQT1iHJ
n0G2ZMknZBou1JkPIiv/ETp/Oja4KcBGDe0Ef53pwZnGUbTA1Y7rDtJuYcLKpVJVoxWnbNqbz6N4
jtNIR83fzgolJeImwqgzR+jKNrkQ6aLrArA5T6C3tNwtyowFhggLQfWFIDIF9ojmM8elr4ofKdlh
LVpv54ICsYxkrPz3M3+Hqu/0hRoJYWEQA3hZ89IlCD9MjQmgz8cx8aO4D2gD0Uq22v0HMQBu0uJs
galEtiyGA8Pt8qbws43TgOHEoo7fDGu7ejVRvKQZzFB/dACLUxJhQ/wfIF3obRUG3qFFgJ4vAYKP
eKPvVOI2TUl/Egns+BhhDLNwQQ1xA7fDoajGaBnxakZWyM9yi0lB/YDwpP9aS4cjaOkLVH2pQgDR
iGwQDn9rvIJsIiYSF1u/IR91Fnq6iFmwz8QZYkKOiLM2UNClbckwv1CeC1Vd9QLoWuPyw52NL1hD
H7rdhh+1n5H4BmakKUDAGsH9exux6ZyQdx4bSZRWXEGZj0WDzmLaTJpXjfCHsh4VO9G9lLOtvQAu
YhtnrntI8GSXdK5i8Ll6AOJEQ9IttATjx3g6JX+FVhtQveatJ7Z8Ks0DtjoalxWC38LXbE+LzmX5
dgbOAZsKBLSLkF5qqg9uNLhjBffwcsxbEh1p2qCJ1dOLDAdBBRpgn+hvT+C1hkf/YbtEmXUX136i
1yq0aMNLkh5qHz5rE84TuYFmVQRKnZqbshQziVzgl34iO5yfO6CQqS7B/ndmiQR6ohRuNaduAL1l
TuVx9UYgfuakDsS+TdZRs2vADVTrdK6YXWeON2brW467oh/A5hu6DjhNXgCsnN7M8aPVMec0HldQ
TQ/KdwprrcMiZAOH2FI0RHkFv7hcEHQ6kjDvh2oSQhGCuDGioORC6XYjEKwQujOr5VHQ5wHUQDjW
G+rmEd/PBwARYQ0xWdZoQSH2fdxsc0uBkxo3ibreOnTHBczaFh9ffXLtcFPzOT0APTvxoiJI1MUR
dGiyg6ndoIAqYmNZzWPJSmN24x3knAv0z1EU5zt6AO5YCyXf63AssIzQujwab8rU7Fx0dpr5WN3d
4wYFem1Ybnvq+VnS86Cw66bwvnLg3JlK9JF61QePbR3EydqbctO/Y/kCw/NEDUtvrnqMhpbgvA64
GDZ1BjONXaY+gp16EtQUT+CKoDO7RPwhM+GvtGwttUBmgn/PEbRu4dx2W7lY9uQTIYanXfKYV0Ot
u6yhZkqnIqe3k/hAYKjycJqVTnXGBMEbGKZgg/Sh4r+ieNv/y8o5kHZL2KUI3Gw4+T5twfGS2N92
/LVY8SKGRg2VptdGVmwiz9NMGMlbxWLh3Z0z2fwjPW51VQLrgy2k9LxvxEmAuMXAKDM/VohpIJgJ
tE4LZbvonmRpelDMrf99lgfNOfBP3kPvcbVuaGu8yoKGUrD/iHH32C2aSuEqWnNSEZOy7aQ2ssR5
hH3U7YUFeY9hF0oPUxem8G05e623YFzt0rdKeqqFYEWDO3H24Z1Q1AOctqwG5PVKSZ/D0YKp4A0/
VPEZGGe62gElBdQcGObUv5MZvius+Hu51WTyAYAOfZTMsWoVwe/tF1SE0bMizJruswb/bH3zFrfy
ei5Aq0K1CeU1d5+MF288R1YLg4T3W5t4Gc1CpkON5Vn1qtRh5iRISIOrMrqyEFW8LOCke89RjLtV
XI9CWmbhVUcsW94h1sleYKmrhePU8ZdriYh0pCO80SAYIUCc6+ByVAgdSnD9Ctw6jBeN23zTCvU9
pNZDfNBsASFLl7mhH1e7VVkI6+3/aZyMWRkDR61nf5bW08JzgXTtPMOxeHaRm4e8lB/aphk6Lhf2
Li3ukru5Uv3DHxACmLh0oeRb6ztC2l91VDwS+yPcnnvEm4NN+ZOBMDG2M00+djM/KJxjZDK19l9H
1nzOmjevFD2xt0wCEeE/Mx+AdaUr8lXIUS4DYoOsErFpcCd2ysWPCeDxSDRAfMwmXiPg7taatlzn
J8jbcb7kzYoMPT9KDVAkRG2quqBPdTVzlhHW5jQc502UymyC/0iyAdmUTO4hd3W7l+BkadYMzq2J
SmH36V9deJ4dWEsOwKjspNvayL8IYvoF3Jcb4RU/15q4CM5bcp78nl4cf0Hq5tZbKkIoILM/aXB5
yAaTNZHb3C0Gw1zhWQ/xBsoebpKeHqud2Docy2NkXcxBH8+7eu8SdDzDQ/ht5qaqdJsgkIp38uQ6
Ijr5Po0vknHwlYirN/HfHwbdtInT16QsECSvdFqnNYXb3VScYjDfxIVxjxRP3rFEYu82HsPxLghK
CB6Im7qxGLWzjdDmdlQEr7n1YbLtgyEF1MdtRoInGZ/wxLIQb6n6f/Roho6LSBNabsDdlmaBRZdb
iwvP/S5lWXm6KIDwjqBEvGyCzsxL2yTJOGBqH4m/ghnxG6KJ/hZMO6+J+WVFIxWh+b2aE3v0yL3T
J6U1GecI0gvc66REYGHKRXAfZSu06iQWVxWwGu1ynQ6WEPrlcGkFU9oH/ltOmet+1nzOoWD8pDuj
4S2gFt5Xty47ovNXC7UN7SXFQnkIllD3n6SVvnhEBEUoFaabJIfKkl1h4fD2TEtwsm+G4+wONEk/
+zy0LuPr2A9vYY4Mij6HWHvB3V43nhAgovZDEzXr/T5YOFdHSYjQ7sZythf0u81yFwnEutLpKxGK
ii0Gs78Gf4cccOfcZeeFLoea52xuTTfhvb8NVcxHnoh5uvmhWhcvIQPs1qPoUmwJwMn65VIzwpc9
adsXtZDx9KUhH5schISz8EX4tbRQkaeGCcVOJ4LajJWLbEoSB1yTGxmq17HxI00QJaEbF2jpcU3c
17TzzI+dy1KMqSX52/ovoW69lteWAuhaTZyZ/nGbGw4Pbs+6gji3bR0KyEviuk1r4fiIO77EeNJg
CEpni0sec9bt5jBmxcEDYAvRaK+tB8eDte76mO5DlyP/8E6I5fyCiMnGxozQrz0u3luAyYhXqUFi
aKx00ySYX5daHvw2JVNtq4alLfWHYJ3oH4SZXSVgsEC+rocbdncYALkVYaqA91CtxxwlWp1kL6/R
z4zg0fMgi/ospUhguWyLOIU0eP9+1oInXcK5fCGCpf0plX2ifGq1VEAtX+eK0EvdTKo1t5vBuLWA
0WEN7eXVK3tSVH9KE9mqbFVXMGXVdcxGny8mp2HW2uL7UCq7+W4u4XJo/nHH9zvyVPt3X19YpnWs
daG3Wws9n14YKbjk8Ck5ctY92DRYGOM0SNnpxGxCEGgdANIgtHIm8C1ohaOy4Vpw2gkdKCwpngQB
uvtH79BuYeFaSmYdc1aoGsneEQhmtFCBmNeuV+XknAl8x8Z33JXPe73MsN5heZh3xwDmJdkME9tR
kNCO4tT5TASQ7oANi2lOWyKvLEVLoc6XyWM4JwmY+CFck+FLn8pmuZ1Uu7aMGHXvihHsWtRM2Znr
Whk0DUjZFmQ5fxsVdGSKFlE1hIViVUstQW73xxnjTs+ZcrbK2PLadW1UlRJCIJuIX/QAATnAcIrx
rACkF5AuiA2jMObksircWedzSH5Vrn/ieS67SKDuu02mfSu4tCCF9VZjejx28FG2TiDZZY0JvNKg
7O6ysxbzcQo+T2KQOKNayyAQyOgrfJZJ5HKXnZ1LPfN5j+nU/OsQeEeekIp5UOLbdFxtStt0ZYRN
Y1yNeUbdGRbn3d/roBL7IaIj3QP+EQEyFqhMfnKCpW0nQMEVvUQXt9IueuvQS0krBxLg3iVCaVpK
Q5b+dLdn96+N48qb2nkJ+zJiVbkX9/CEmR5fdtVW4ruFGUc2VFhXkj191IzAkabcqZjZNsk+jW7p
oJPSHIIqgUkjDsnmgWOr01Fyxvf0plaf6ctxx57eqZ7jd2YUowIsZzBlcUFxBAr4FRadCf3M6TLW
4ndPJpJuFAbFrEF3BeQAAKl/NxJWsW3yg9k2z49DKGpI8sXVCKlJkIf1OgI/WUqz3IQvhQMYmbHj
hG+dyPi+qOmhRTFSybEjuy5VD02Z8XNDG1h5OPXRq4f4ocT9wDXd/IH79KlKtVahRYD2fzwIvdiH
pb2V/BoiRrjii/4f/Wh8XU9XDf8N20MQPaqjW6IycrEyFH6B01bsZWMGsQCM8lWlPNd8RX+dhWHo
URrM9VqkTX3nhkt9YwUbtR2IfBo0A+17dFOWnKs87M0UtWp2X7Fl0Z72dbV/ScpNWYnt3Sqda0S3
W8oVT+HteqodSzk5Sew18aQ8FbITWZE4Fjk4Bcl/0fHcR3jTrK09yf5NcWRbFTWcPqnUuIvNkpv9
91s8f5XeLE17v7bM02KkS/vtc4V0rXf564i96n5YhQxEFXBpwQtiiF4yQ14dXFwgNLlpj8rfwVdY
5/i8x3KbH2OxFLYbvbP3BhI46T2++bmbmMX2GdY3ZJ//BWSgAtkcFYHrNys4qt0FmH4tWy/CMi4v
DF8L/QH/QHRsyEchViEn1oCZRAemQVIAB0+OFdIOVEa+LESKFXiagMPvcj+Y3Y1OiXAyUzjfoOeY
XG8MIjyYpcWDPD02sxPEa7z0AMDNOCLFtACiR4C7lOrLLIkzTHINs2e7yYL+6MIIxvIG1OdBIqmu
ZH6xpSDC8Rf65t15mno+x2qhyCIlRN+JiwlO3isUxtkmUQ2aqSmgfUx4JGwTbwZ2YNhgCpROuXbX
0pQW4YTP9ab6eRQdWzm5tqMyZJ+vhctq7Exz5OhWjQ28T5Hkd3ejCtXkvoOn1cv/zjq+JnpktoJQ
KJ92bRrxEIfEjz2akrbwgbOeoAcJy2E2nG9ggQxpYi+EmRfxJ0BQfS7eseVm7DO5MhuSQd6Y90y/
uvAvQTPjbXio5c2bh/YUn7t87xVgbljyDCLl4W7QIYhQ/uW1sk1gWcXMaHdhZnT7qnEmtiLa7z2q
KrIHTA6Vv9iNtLltCq0iIeCFk4zpR4RyREoozEEkHKK5llz7a1Xb5eup3Mi16+KzfTB4Vi37nsM+
cHRxv9MSs4JMMrDumqj7YKiPikj1PfJNFzSxEL6IMQisiiZsHQbc/DzcSfrQbUS16GKCU4AYnRhJ
ipgjfH7etY75vOT+OEgm+QrDkahWpQGmCjemLQTIGx1ZMkCO+nwj7co+muCBZ0LVzKB1nlP23tow
oq3Qici4fcr2vpZ/OqY7Jz5Ju5PAc1EvK71DTKSWfDFTNaKLsat/0zh/PaBSwB+Whl0a7krcYdWx
bwrBPnc6a4yIy+dMn6z3pLQJmxEG61sQpXVQDISkSRy4BTwv7EldOi92vQszOt8sROkCUxJH+xfZ
3DHLs97JMrSflgrDpzw2g+7EO0V2rGbpyvNyEQAish2rcAQnLUfjTIubCoRJ4cs3yAT8COgQTP61
uOOuCfzP8BlCtXlVs2BvbkZmwpzpf3W/u7rAHosvMU7iwiXDDTACuEPUArVAQ05QsHTL5mFuVh4+
R8h+weJaDmxHD6PwgCty
`pragma protect end_protected
