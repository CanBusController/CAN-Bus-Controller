-- CAN_CONTROLLER_tb.vhd

-- Generated using ACDS version 13.1 162 at 2016.12.22.17:16:27

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity CAN_CONTROLLER_tb is
end entity CAN_CONTROLLER_tb;

architecture rtl of CAN_CONTROLLER_tb is
	component CAN_CONTROLLER is
		port (
			clk_clk                : in  std_logic := 'X'; -- clk
			resetn_reset_n         : in  std_logic := 'X'; -- reset_n
			conduit_end_rx_i       : in  std_logic := 'X'; -- rx_i
			conduit_end_tx_o       : out std_logic;        -- tx_o
			conduit_end_bus_off_on : out std_logic;        -- bus_off_on
			conduit_end_irq_on     : out std_logic;        -- irq_on
			conduit_end_clkout_o   : out std_logic         -- clkout_o
		);
	end component CAN_CONTROLLER;

	component altera_avalon_clock_source is
		generic (
			CLOCK_RATE : positive := 10;
			CLOCK_UNIT : positive := 1000000
		);
		port (
			clk : out std_logic   -- clk
		);
	end component altera_avalon_clock_source;

	component altera_avalon_reset_source is
		generic (
			ASSERT_HIGH_RESET    : integer := 1;
			INITIAL_RESET_CYCLES : integer := 0
		);
		port (
			reset : out std_logic;        -- reset_n
			clk   : in  std_logic := 'X'  -- clk
		);
	end component altera_avalon_reset_source;

	component altera_conduit_bfm is
		port (
			sig_rx_i       : out std_logic_vector(0 downto 0);                    -- rx_i
			sig_tx_o       : in  std_logic_vector(0 downto 0) := (others => 'X'); -- tx_o
			sig_bus_off_on : in  std_logic_vector(0 downto 0) := (others => 'X'); -- bus_off_on
			sig_irq_on     : in  std_logic_vector(0 downto 0) := (others => 'X'); -- irq_on
			sig_clkout_o   : in  std_logic_vector(0 downto 0) := (others => 'X')  -- clkout_o
		);
	end component altera_conduit_bfm;

	signal can_controller_inst_clk_bfm_clk_clk              : std_logic;                    -- CAN_CONTROLLER_inst_clk_bfm:clk -> [CAN_CONTROLLER_inst:clk_clk, CAN_CONTROLLER_inst_resetn_bfm:clk]
	signal can_controller_inst_resetn_bfm_reset_reset       : std_logic;                    -- CAN_CONTROLLER_inst_resetn_bfm:reset -> CAN_CONTROLLER_inst:resetn_reset_n
	signal can_controller_inst_conduit_end_bfm_conduit_rx_i : std_logic_vector(0 downto 0); -- CAN_CONTROLLER_inst_conduit_end_bfm:sig_rx_i -> CAN_CONTROLLER_inst:conduit_end_rx_i
	signal can_controller_inst_conduit_end_clkout_o         : std_logic;                    -- CAN_CONTROLLER_inst:conduit_end_clkout_o -> CAN_CONTROLLER_inst_conduit_end_bfm:sig_clkout_o
	signal can_controller_inst_conduit_end_bus_off_on       : std_logic;                    -- CAN_CONTROLLER_inst:conduit_end_bus_off_on -> CAN_CONTROLLER_inst_conduit_end_bfm:sig_bus_off_on
	signal can_controller_inst_conduit_end_tx_o             : std_logic;                    -- CAN_CONTROLLER_inst:conduit_end_tx_o -> CAN_CONTROLLER_inst_conduit_end_bfm:sig_tx_o
	signal can_controller_inst_conduit_end_irq_on           : std_logic;                    -- CAN_CONTROLLER_inst:conduit_end_irq_on -> CAN_CONTROLLER_inst_conduit_end_bfm:sig_irq_on

begin

	can_controller_inst : component CAN_CONTROLLER
		port map (
			clk_clk                => can_controller_inst_clk_bfm_clk_clk,                 --         clk.clk
			resetn_reset_n         => can_controller_inst_resetn_bfm_reset_reset,          --      resetn.reset_n
			conduit_end_rx_i       => can_controller_inst_conduit_end_bfm_conduit_rx_i(0), -- conduit_end.rx_i
			conduit_end_tx_o       => can_controller_inst_conduit_end_tx_o,                --            .tx_o
			conduit_end_bus_off_on => can_controller_inst_conduit_end_bus_off_on,          --            .bus_off_on
			conduit_end_irq_on     => can_controller_inst_conduit_end_irq_on,              --            .irq_on
			conduit_end_clkout_o   => can_controller_inst_conduit_end_clkout_o             --            .clkout_o
		);

	can_controller_inst_clk_bfm : component altera_avalon_clock_source
		generic map (
			CLOCK_RATE => 50000000,
			CLOCK_UNIT => 1
		)
		port map (
			clk => can_controller_inst_clk_bfm_clk_clk  -- clk.clk
		);

	can_controller_inst_resetn_bfm : component altera_avalon_reset_source
		generic map (
			ASSERT_HIGH_RESET    => 0,
			INITIAL_RESET_CYCLES => 50
		)
		port map (
			reset => can_controller_inst_resetn_bfm_reset_reset, -- reset.reset_n
			clk   => can_controller_inst_clk_bfm_clk_clk         --   clk.clk
		);

	can_controller_inst_conduit_end_bfm : component altera_conduit_bfm
		port map (
			sig_rx_i          => can_controller_inst_conduit_end_bfm_conduit_rx_i, -- conduit.rx_i
			sig_tx_o(0)       => can_controller_inst_conduit_end_tx_o,             --        .tx_o
			sig_bus_off_on(0) => can_controller_inst_conduit_end_bus_off_on,       --        .bus_off_on
			sig_irq_on(0)     => can_controller_inst_conduit_end_irq_on,           --        .irq_on
			sig_clkout_o(0)   => can_controller_inst_conduit_end_clkout_o          --        .clkout_o
		);

end architecture rtl; -- of CAN_CONTROLLER_tb
