// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:39:01 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
mXTHl0Jxj3aV1EpM/QFTZd3zoe3XlDRRdnaEXaTe/RrRujMClsqUQvTuuMaToaAj
V6msLESqrFurb/E8Sn/Y+A6OLFcn86NTElpA5AeIY2QmXSqE0hdDPKLeaAestClH
qF8delKsgN6/wCke7iN002pSKXer2qd1Z9nKPwYWrXA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 14016)
u8RyPZNqvviST6ytjkzS7Yo/QgHWody4dZKOFBfaIKhbioXvmN9PTM2pO8TQ0Pzi
aGj3iZpO5+MT4xIPPJ+BsMhqeHKqILVMrHwTkbctnYWB6qkhSBaVXsRrM0Yl7inu
SKpvPP2X4bduQEmcrjS3znmBuF+VliUKAl/6xB84CWO7QyKuNDpqnaR1tKv71r50
6EDD48MZg8S9VahyxXemz+BF6NLRTupqI8wGblK1KlR8xNIzhoUAsq70optRHhN1
lwfzzIaM/b0F3PF3BnPz9H1TB7UEjm+htwCLe8h008aDvpdGVpNV4Xd7kzFE72q8
kR5h8XlyIG7G2pM9Zq8mw1jbMNNiwiISGzWl279wSxZOXoVi9Hb/iczy/v844T6w
SYTX1qdOEbCmqFVc0ur82jS9eA/jg6wau4r+zuRkUFcTSuz9udfB3GOYNTVO/Rh+
vrh6Iv5qPRpEk3HtKAm8i5FT7Jj9RFl6L9BmeF3+plgXyV76OJw5nkAxRWofZcnb
lW786JuMSJMssEKUatkqp3SIXzIT59+xJVbSNnuc50ER+msc9kv5xST4lJRV+zUB
f/hWshHrx1Hw7PRVE9CMCQZt9URuJoACtRValhDwyOo5P++eqSIzzbjiLWay2SKt
zE7aljlcuBu7oiLs5iui5k2O78m90MC0VS8YPNQGEQ5oEnp6kYuTKTdJ9Z76pCaN
MHIUWt6S6ytJEyfRUf11a+HeiLkq4YgADa8e4xd0FoZLWzQsg0qHzRFl7eGqO1Qg
N76O7lRq29vNFQ8P6grvDvKlQzNZrOVP75x0az8R9C/7x0e1t5LshF7t8vMbR3Uj
vsAMizmHXeyZvBk4boggXkv0ie0fk2LlY7jzV3uVFbFvVfBNz4CAboUYWsvDFin8
gCMWq7nG5UoP9sUNb5tRB1PCvbVZG/AW2oNZ2vYrwG1JFqUam006kcTLd4JfWfn+
7lIX9JK7+r4Jf9o9Ick7nNKrU650egygaKh2SF4ZcsDPFyRQgDH/I08sUTuscVGz
vDSslFb49XxQz4DJiQjAfR7tHXfr+FqFIzoV1GWtCP7/76uwQD6tluSjCAWK11Dn
MbHxI7XLxNwtjVc2EVBXvETabWFoWY3DdRUuz1X/BL6DJ4DAk9/i3YbO7bjirTPe
ObbjY+oXU6BOViw9pvVCaeZZQPuwGL/+BrNEex6eg6e1xS2dkGXrqlZHKVtiHF9Y
UstLO5bbpXfcrac+dg+PfkmNC698Ifyr17k61DXWrNegTUlPhWDrZkx7us2G/AqI
v/GuOTRHGkVvIqg7bhf+X/LAR2dxaZrD+1zDByottSG3rwSBcAM4J1C8ZJl3If19
4PrGex4dKVzETZNE/NBfKkQr0c64kNncNDLIWPSElC8klcjPfEdoQbtd+OyzyJ71
am2LmdAf+YoTX7m9324CPR0hQdwxBya146AxOj5CuAHEIShb5o3iH2DsKWSTIcNy
pMXqMdEKt8Xw1i8dxiRZp4av52Q3VemNDx5RsKvf+C8ZK3ri5YelzVZal7p5JpPc
tC88PEqjKjRXxKJYCuJgWinS/zgepY3Aj11ioERxzbJcrf8/KveUnMjq+W0NM87H
vLcexTpnHI3z0j7OVObCcrelItd/b8TSdF1wO5qV2CDvyxvvaRo86cfbgpbKYs+l
DczLSe0ZYw4HYQBAcLFLlEvhGSFqKf+89p24OJjWj72O+5mLh5hNSJniAASitjWr
5TBsn1Ebm3EaGX6keCRbNIIOLTLCrCADHUOIFyO/f6wBO/XBSGBPnklrNVM0OgDm
+2gXev0g13ieCH88/s+QiFrT6R3D5Bwx624FMjxwLQDLuPS+CdkZwZOUbIgn6E/v
icDcZRozMwYC4KM7VKAe4QWgCI8WmpD1j17YsBhA2zTxxFwnQ8FqqNaBBydp9DkV
9R4uhXEap9mCTpHA2xFf1ePk1XwCsPIHWV2pUzq8DEqxmVYwSngaEKuGpMFWVKww
dfr9YHtX03LdeZMCIVuaxhinHJhiOxvuVvXT6p11gnPvdOfb+yXEXTWj+/rduD0P
jB15KYugGsprpy4DPvqJjM+YMs6UFfIWH545t1KqE4/PKfNNIfrhyt25hjWgZXaM
s4Lzyl7NTPPqyz5OXOOfqwJy/JU22mb8bNd+hpyhIbhGiyC1JvokQb+ed2mI+Aj/
i00jNL3G6zkYhsByOVCGpm2bbDWvbhxTjhIko42N0Iv05Y+lJzw+o5T+Ya/DScUY
tdCmjQB7fQrvdhHi+0C5PkPcv/DBJTLMAJue7W86UKFGIH48yit58zV0OMC5jOhx
c683IobCTwkrq8D/Jc/E/RsBsGQGUSv3qn7HCIgktFdiam91wMSID2PI41A4lw5W
Bka5fdXsEyxLVccEAuPJSwGXlX1cmah8X/qL9ojrFpTuFLF5jI9oRbqqm/gWN0OS
yyRomvmHJCvIa42zJdn/5y0xivfkpjYAC/7IMjuEk+wsqKMHa0oV5L/Ax4hkbOsx
gioK9QKojiKG1GnJoeRRg922AFZdMyLr3jaLzOQ8Y0k7V8XJ5maKui+9E2OtSvIR
uTecu9ojKMUpJLrIOn2i9xpygKefJnqPqmI2rs+peifjnYAEvJcYxApn+xmS6Ua9
M1Z/qbCrflNXhLzKb6Ydd+Fknz8XL5tqxzsy3otgZLgbnkOHt3IEsBEdPVpDoBZu
JGyBdbQSkYWPWs8/Kd9Lw3rj9BqyFgmETseaCEVAtkVNNEeDj7HBeH9MYqJepEb1
WeJfxqwcX/mXipacvJYAiBbVCMX6fA8+JZdRzp4+K6rX6sJTdkirkpWuuQMO2sUN
GO8A+EXrneQo07blyvUD39Ozy/epO1ptSi1esrHbNgpTFHhEtIRFO4TxthSmGTya
ZbRHBtu8ynwnkkr3c2oqiCzOQmjUlsobxcpwfabZYEbVvvqDiQ6L9PVmrS+JA20m
RO1x2gO7Q/0TdsDFMtRS9q6J9qQcxeZRpmaIHBWXk/bO46VxyPgGgk6knQfbqYNk
oj8rB6aeIn3AHSFmN3h0NXHvnZaFOW760iZ9xRD05HMXC2wG13fPJlMXjcQyP+XN
THxFxftCiWC3Nev0aSA68/TJpDvSTWHjla1Ie3Xpbty8Bb4sMlaUV0GdExUk5pmm
Oz2YZxHPc7PJVaUTm8/4hOZkEd3klqNCgJM5kAhskEfqVn9+RqLS3wA2DuY8B6Q/
EcPVfaezL74L4QRlFqZTfuoiN+vKB83IpER4oC+APZ4Rk3vKHcGR6AP8VMY+iuKs
dZHwKxPvKuS8t77vDMrlbXgwEWR7SEfErt9Tkg++7hqc5/84IY85Yx3xgzoJJalh
SjNqc5juX1nd4ofvSBmjTtdembBp7ntwvXT44GpveuspB2cD5m67Xpv/Dbv5WwzZ
uB2271VPLnGs5833txrRq1WzqjnJrYUKM3MgABt6h9FNcjiLXlqt/dOoH5ArkWI5
0AA/1aKYaYXul3BWkvPKjOipEmoBnjAIgoH4EX0vMW4SHVVsRGslhTNrCrqS6XCI
xncEVWm0447HiqzEyg6T8RGtsZO3wjS+ziHK+roVm4SDWBdckHXqhC5rgl8uE2tc
9pPnpwXUBO83LufQV8ThbxmfLBa4u1wqylZkQJWAMS1U993WOzpfLujfLooJIuA5
cZl6cxS3ic/mbhPkmikHoTEr2nKel9VjSb+Y1RoK0hE4z5FJv+VXrYr9KcTsciXy
eAfgXoBFQjvFm49zwREBh9qPRQrsMUzv9/KQuK87Qgpq3byS7IrEAPD3UiURTtYJ
RZaMuhaZGjF/Ot6npLTk9UboINdbQnASYpYF7XLdfxuYmnUMV0gd03xqs463uoRA
GxVG+uWGfSpMK/W2bGfFVABN7o1M8WtXnv8mykIvD+xwhXVyGFEuU0eP8bhqreH4
XojJ3ffsvpp2ARDVrNB1Mmu1SosWV+qdNUiU3j/S1s4ueP46N3bm63D+eJG8qFv3
lVWGcT48pRPVlMOOoHcUbjwXoo9xgpWYfkvkhY6dg5JqWLmuERbhHMaewWnoJ46F
n8cESyLMPRyOvmnVBObRyIqhMQd+XStP4biHFc19NoflAUiBv55mbC3T5IRP27SO
OUxEISDEWxouyE/T9weaSRfEqzr6eHn9j7sLwRbe+SBSRIIzwfN1irQ1qRPr82oZ
+9Pzkvf1DzFHefTblmQ5W6zh5mV3WRcS2pYbj/TFGKlAnrymSS8lDBLesWsl4Zn2
so8JwNp3f0WHVHdn3V2ASm6jel365PSh/TQCExA2ymFy6mL06obLBiGzwPkOdmI7
1PUEuuLOnv+9GTMt1ol2DhXaabaP4mkOr6kUuo/6Yt4/cPNS5cUUQUDHTOFBLR9k
XaG/N1lBLisRxeJ2AJaBNk49bDq2BBd3asetX0CMyU4b4Ub+NVjesKrrNA2z9ZU0
peS6kU+RdHfc4XmCEnnGq4h+z3B45EgpmxthzQ++jLIB5EzFS9fyjfJK7E3XKJqv
WSovOGV4w30Gp60Vt5KsZCt3I0dANb300m5fLKkVcu5HqbQjzwPWc4X81yHrvyPv
mk5PV4IQu6NiSO3fHOCj1tbIrCtwVUMur4WKj2gTWJV8cAsKwiWko7vtefT2hGXf
HWSW12tUrwBWhFXLeYY5ndsvJqILrB6fF1n0ctaMfLwwc1M0lRhYyxx/XiHnkWfr
kIPZAOQPoRZ4hvUAQ3HjaE1oAsyUqCp67zqjA6/VjMS4LqoW7DAQrxut0Rcu6705
wQTVaBO4AN45H7w75XADYK1+2QgFccny6BoENW8/3H41eV5/V1sxXyAYl28hteeq
t78c84rY5qguWjCdH1Ma2dZnfJg7eqOTWYTh5B/E3ZD3zcd7IFG5hdlrAUxvtbkU
c1xiK0a2zB+Q9ENdBLL9T+fPAIUtk9SCeILKm1tc5kZ+l2oRHC1rb2DbINJASeEr
PZ78tQfmYbCuc+FjTu5bg/Go/qhLBs6qbr2mekTVNbjaCWXKWHzZor1HF9qgul9H
E+SGMGgEW7NYKENWONX016r+bi9rAYq0CYLnYUqWpS1G+t0GQYWhzW5oIHIrcvwy
XvO2P34gYa+Xs/KppqZeUzHznOx+YCLqQGm2/Tco7GxwvQjYCAiRw0ghQe3Sl379
sGEol9r8BrTCY43lEb3Xow8seyFV9EZ6u10JstByxm5wLPEgyMOuU7+FPfdlR2J6
Z/xRQYp7IQ4Tw+j3Y2FhfwtCdJvHMfOAHkfYIgON3b9eOGeXD1JQCbvqHTvz7Vic
1Of4X7KgY4jv+3x4V8IjTU2CN+komX7hX5U824kvp/9G5o8SvF5ibqWOKLPTZQDY
N/UJjwFY9+FmdMIGhOvPaaLRnZP/KviyZYN9hr5forI0byeVAIaXxiCHYy4ni/IW
T0BMubgeia6SD2xFDLromlhUY0rR6WXgjaZskzTxp5OzKRVAiCmG0CUfAQjaRViA
m2bIqFKtDP8Dwhhf89M8ifxiu8tcfdbV9TQUWx+K/a++vC2vq1jzwnpohlBAknZY
b6NaHndocYkwRtIfpM2tdIHMkOrmh0nPHuD/fWzLu5nKjGJLxvZxEXShn3OiZPKh
tvle8FHITs4qjFoUmeFG832AKg1r0NUN1os/jP2Q2v73D36nUy0a8LMEAXdQ7E9O
hdYnriVycW+UL7o7A+lvaHeeXh4U/q6eARMo8ejrvKmSOG8DvfoXEXQbQWVwH5XU
wLZ/WVnclFjW5zOnrT7WwH1QUy8bR25mQgiTXS+r6bWQqNRhTEccJklKYxFZoDZI
R6np2NY7NHtv4edmxh9xDDJfBHg4QP45XFVDfdsG1X2d0NeKflrxNaGSWYJivKDo
bLGFFUnhrwKGRtg6LKKNMPDQfMXrFIn0Mbl3MQfkcNxLwCAlWahZMySE9QVg/Bhc
oob8VQKxJZ+qx0TLnOBno6/5bk4qwsWy0srEQX5f9XN4Gxz7p1yOZbO1I7/0dKGy
lYeilWaNxhB7rt1Kik7/QfuFNcjosMGuI19MbwUyVXgsOtmSWcKNNS/cQYZneTWD
bKCM6GSLlimEa9l5Oc+ptLM7RYdVSBX34WNTD5q7tJ7K9n5pOj6xoLNfUivlwHLX
EpDxv7/jjH/W4hvNFR/bg0KRoiJAOCDTxHuFRiwfBOQwSSNAH2yy4I6RN1JocD+Q
LhPLVhTZF1lYEwwN6lkTaAtQpOFa9OKUxuXMtKWYO/MW9C3cHG3rb3ayBVCTpjzy
Bz9bjaCsYhfEJ+NODbB4K3r60u+2NJuPceNz/idvZ2Os6MZhkIaRUEhlf+fnfQ9x
C1oarAABcdvS8xg3AnL6+KfiiHROpY9uD5/8h/Fub13t1zUkCS8NZCEpNTTuSjB6
gJNg6kqL3NM47MWBn+6M6F7IwS/lW1LDgqbvZprclFVgOohOlDb/1v2EtqA/0UA8
BOC3Bdv2KC+vUQ6t9m7mPMyO9MKFqEqViskWt84DAjRzKyapxzTQL+zkuHisZ3Tg
kTLdsB1jRXCFfnZls+KaX+ESwAQLVn6sHz5DwQbYMWWrdgBmqzI5E14GzUBnaDFk
64CUIv/Xtl1dE+yEnsHNLmS7qQqWiWDdw/RSMaYQMRxAWggbpDDbci83JgPCh/Wu
HltTpTmu4Ilc5qY1lHcVry2B2J1eiCTYU4fuKy+7c2S1i55bnH9wapgVxLXJi+eD
b+kPZPqHw81RjZvZYMc1vTEyn4u91dc0MrKGOLvL3flYw8ZdzCJXTcmvI1iMJoQw
DqUcbzkPnIMKQujeNAaDxpXsF6ZePGIiSWI5r3Iyi6sX6t3M8J/RbQdhjuQ4bhHv
7MCVI/s/A+6zae9neVCiRs7zlw3HwPfLuFFrBPTkO1G62ZIvT0EEwMGd2cbia+De
HU/1HFYOE+cVtaLlrm0l9PR0xUbK7jvWT73DYSUPguGV4RKc6Pbq6Sx+lyaHzYg9
sNMR9sY8lDdd6pFq6q1TiuWfKIbLi+otPETn+YNLqDsEZQpbN9QmeKHffCMYrcCL
mQjAY/kTHZPF5G84B6XlcInTL3ZoMrKAHQD0EqIQ0pXzPAKzQz/pcUw5vKx06In3
cw71MI6n0jV2tbd/kbUq8iGn+c3PvnlACVtH9G1OsjvVyQ0f7Cu+M5/RjdZO40D/
/PPUYDelA+4CA+Eto32rilg6k5n5SbtBOQyuD4+XUMrJFLjw12lJfRkTQ7gyOS/q
zENGb2zA02E1rQ0OMpo1lgfWQ/vPj306V+vGyFwkkBIMDIzSQgRZqhI0ONvEuqIq
Z9iBqA2MiyotmfcgCzoRhIoVMTwqiRTm1nmeMy6p8Zg1MM6lWB4+FAgk5a33idv9
0hsEEJ6KfD5IJfhZvM+lkw/rj91wGoWKcTUfAQQY9ufB2W9qT1HqMYeNyhfjipYQ
BdyBSGm5XlZIGlxLbNBXwAZ62EmtsmiVkl23PSolx99P6z+OoJTNtYsFIjAIo0LM
S2/W1M1fZ2PK0ztL0ny2pl9YeFNKmmJBOTBVxRUi45XS+tMT0HwJbQaUP7kxFDoK
HYmoTJNdtAYHvNpE7vElNU/2kmU2LALcxaoLM9jfYU+UuryJouf6IPyxjtaMS4y5
n/MTsFkuR8STgQLDgInDeVS7dG6WZJkPV4mmYNWamheFQ+9DpIeCQnLrkAR/0FwF
tWTtGdTBfGrjFfWYDo0Ry46Zs4KQ96X/VqaB5rik3hM+yYUYXd4BeuPuYV5Hka1w
fsJaTb+LXGI5Az78O2pxea6j6+HNaGeFVP2inVqu4cZ+CgTvszQws1pZvvIOS+N2
XIu7YWlND053GnDmkSbPZJ+usRbEHx3g6CxHXOooc+ogdG9fOmot/KJUu3d6HSk9
GNfhcEbslhCSBHXqOg/NmicKQmHa2dQn0NjVFwYVsLsdqc/VK5N/y5bPL//lckLA
jgsiKRzzQcjC3SWgQespeQPxzkcGYR1+NnCoYjTWh28hugSdULjgy0KQwa88TrcR
6TkuvmB43WC1BBhnexc8vR5Rw8HRYXRvbuqZkuvIYdWkwlKMb4xZg7m82Q9ISsTs
iJrcreAsB2Rp7CdxqTnyMmQPkzqvzq4OTzFICUJ9kwIIrqzXS/NV3jzZ0+b8RXN9
wnXxutwTHSwq8ndI6yvQp4n9PDzrvr/OKNYwRvc7pOfSkx6r9Bj5lXQ0xIwq/i3z
0/OJFWfMIcBgnHqABEqIhuqEJw/l5fxw5i7/lSloLWHKFDmM6GuSSFDiY/rX6BRJ
cd+oMX+NfeTDzly1NdTlkW5QYbi0BmWyvAshEYtPC++uYBCuxLMZkd8ywiQEoNyO
TYba0IXTHWnvqoV/oHdSBGHx6enI3vx+A38UEiKFervhRZbznS0Uj6esVctKCoCf
yhRhbXpswy/Oe0almhmO+z7Ep0uKGfj9j1tFyr7SR/yRMx9155iHJ45S76boRcCw
ur/GPBnzLu/WeEWA+qYY1+A7M9Z1ulNM0E809u2CcRsbUc3Hz01F6+rTddGdld22
UyrOm1aWzog2HA30u9QkheHqs/ld0ZFo/im1XvQIn2Wd9+dl3URkY4fME6TZQTHg
SeHxbSXJx1Pxu03TkBQtM8+/9oC3cTzmSObONccUBYYJGopAnEpRwURZZKxlyhQR
sqy5SHx/R1J6t3G7yler01aG2ofWx/23UsIkr141l96GD585TM6HbIlbECKLmNNT
W6auNL5a1c2886gyvVsUohvCEsYQnIFrsymfpA70gEynC0wlwCA0eHapRnJcP3vx
5mkMVeZTcsNmjSg+KdjwExWXlAY+HRMwQ4pqV7XZsg3FVLB9pajz7v14CqsUlmNC
sLdI42aGswbd+hmdJCUEWTMZOVlfNN89xlK4LnN4D4v9MQrTMlGN/XooaoDY9Mv7
4ukOlt0HtTNck24yp3f2dgnd6hXZCPOtPMyAbmdvOHW3RgENpEBcKs9s+VFuBcEY
RX4ZlOSUvxZ8UO89oFCuXAFRwBJdjdwfIusMIpu/+h1QjJIpDkubmELbniMIqWkJ
CcS53R3KcxTZaQJwvPavC2LB6ew8JDK6s8WYubdHGNZwNt7vLxja1l0VEcDfNjgs
hiISs/3ayRMS8wXu95U3B9ez0kn+8BZ/h5M1eltIekR0RsOqOiU2IkiWTTSUtBZ5
BQBzCv5UG6NyTq51xLi7keyVS+C3cTTXWy3hYB+PxFsVu76AVHh/+dsc9N910VWi
clPSSj3wgfTH+qBRUkjoYhGqk1SrHscGFOy3gsOXcKCIVWegicIHTcsDaa4mamhb
zUvrm76zOnSEyVmXsFQO319YjQLPVAQ1MoFz/BlTBMoECsmM9ETlVizTCdF2FRzW
uwtVlsZkLPeeSYafGT3u7gjHqDMN4G7k6Vhk7xynDWNpkVMPG8Kepkbr5xe8XQQC
3JHTPRP7zC49WOHBGafa0VPLeEhubpGH5RKSZ3oJmGoJ1QHW9NWAG0jAJKQXNH5y
R4AS2idl/BW7PnDmXEPECGFWYdEboSwWeNAHm+SUmB1yWaNgQ+y5fUSCsiN3oJ9E
5UW5Nbd1MQxvy+eU7D/hm1H1WNpC0sEi/HqK4ZHeliH9WoHs4PLsQ/tgGRkTkz11
V3Dl1b6Y10PVOTQj8BrMw3tcEb5eMLDrzZNLa4Vuy+eEIsw38q+5WtB0cUzf472H
ZpAh4MqMJ8V+MTCfDqYYNQQyiW7uiFWJSC93uqSx6DyRbuN7JFTF9c+t57BOV69B
UbaIxnoiZQS+D3B4ynyImCgBBw0peezsPTexezdU70vLUhO3BclLFZjGqtkt8MS2
QFrXX7bb/mSK5N4vCo0sdjA7aUNdPZ4PYGfYdw+RY3csFpnIHbFcqt2i7NTNX9UZ
urZUQL1UQLL7BuFNQQUAUS8INc088pp8zKabEscJX0V0Vr42zTOwl0axM3eosb21
0tZRc7TaGY69m7EN83U20auo+m6Xfdz5p3HwMKvi4CdYN8mbSX1YLEveBZD7tStJ
RvvWaNCqdydvxDkBv+AEbMIT8gWNG/TzazY5B0n8OwUwALGWhI1mdJpzGmJNxkF3
Liuk9MMVAGnvazN/iARE2AtK391FfxxUEMCzab9E9LZmHiAp3wg4w/FMKoChgF0f
MHZa3/70FZUbr2COmUeuSy+2CtBDexK/I8AXbVA1jbVOnoWJt9kxdl6wELf1RAbJ
t4VRSRtuEQ1DkA2/IFVcxjkElbYUiztkZPzJd3MuGr0jJ42DGstQBuqNCH7j6JoK
BcyGWs/lTDk6+4kqmn0KPxAjIZ0HzScEGJ5s2pDFeh9jBbvlBHUssCjxucLdfr6i
vF3Mee+ge/sPkJ3/KKzRESOzVI8b812tHI0vmK+C7rRh5yw61mXVjTcA9bDrsk3P
JYpR6QZzhblrTrCNUHXDWg8FfxuJ0A+TTk11qsS+pUqo3vyCnEAesndBjUHm2XMJ
6y3zOe0jzTNC0a+LQYWjAW8W7KU12T4i0kPl9DXzeaechzFOC68UXlj7ch67msAA
OXqeq0qwg3sb3Hy9SyyYeQYdOmL4dRzHTCnaCze9/qPN5SGO6Xb3hm9aooWum8Pg
UEusmZ10q+1hD9/o++Rv259RfstXFigtiAa2SXMAb9hoBwRQrSJgf8Hf3LieJZ/K
GNzIM/AZ+ahMkQEatfs9MqkaZnU475Lar1WlKhktbpXc9x7/Ut88KRDd9XxQkmya
HjAR+fjnOZlsRRvjCWpCN+Pns9/z2t5TZmE9BQdanMudicpsol9wewH0oEuzG2u4
XxUYJA8GWAQbKU6I1OZAlrbpauBgjgcvjC0MqKyisd3jgksSBYoxx3KnDjlYyI+C
cH6myObBhbW/uRRgpbg8eIpL1N1DKXQvHsxxMEr7m+/OyD+aarLR3kY/vXWdG+Zd
gwkv+GeiLIoaDuGGj4nkmZNZfPbiQbDXLpJxHaW2GweFyFmxZpOFYvkQrzNqmzya
U6P94CTtZ8pMpznokjWmSYmHFsz0H+v/oTjJvvXXthXKuMO07HoDuxjq38vKgg80
UuGDZkZV9ak1tLg+UUFkcLwsVCy+ERKjRMynFihJNa80gtPdvahf8vFlV1HD7cQ6
vjGg9J2lrjlwhOFbj2jYsLfDzkKi68wAWggv7Djrb9k2rVmSDlfMkI4mRRCv7Lii
+tmGUjV1/8axDu5YUlrswhIWkDkSNQr4ZpJnl8WaGV3OnRVyYvAaITl9ewvJhM59
/+h1ScRPCoOWQBFe7tTRwbIJk8vDI0XXe3NDeb6NTqt5zES3n8Sv9kdSHVdWx3Kl
HUKWi1Al/RXV97uB68MBvJK7nmSPyI0j4LSLf8vyrZunkfp6Uzq324bE9yriv7Qr
lTALQy5ckC+S+uCiQd3eGj2liTYsgL703BFA5B+TILW94yXBu5sCsUjgTSCt5vz7
BLhYniKvTumDJcUK0ziS+PV/7XDbw1uRB8CF3ailWBICVHgY9esDBdsf9jY/fAr+
6KGLDY+ba/LMESpAmPtt9CX1GyPnMu6DnDZnHHZAwwN9OaOThWXi2i5YfG0zV72g
cpGWlNMWwqNKji+5fpL4IgwuG97CEJxgEB3NO8/hI66lgjYOOYLUvpbhKA7r7RUj
SBG3G5TbE0zEtBCdy8rebpQXhsWFXFVO2KS3XItt+iDHbg2EZRo9KQ4sCQY28VEC
uWALZ46p6Hq7UB5nEFym0hiN3yaPD8l4i5/c7F9aPaHBrGqvop9X631ja5YUYcKd
VENcdzC4svd0eD0nqj8W/Wv4IDe7vL4zmcoJ+vhBYn38fx2SfoD05dUFNN0ynZ+F
VchsL0SPlMSWWXNyBQ7+5dMZV9qENAAE356PMGkL8YqoFrF8LFgyPJJC8ypNh7Oz
V7jlw/g07EP78FUy5PUvKYTJVxln7vwno4GzQjeoo1GPJSLVe5k9hqZ344fpL0O+
7ePhan6RLCvCgdBvhwp2TG5sz5ScYaJ5GYrK42/s3JbNDuCDJvYniQ05Yd0GhTfR
dGQZ+3sEPA8ACxAAzvRiw7XaSlnN2YCsvLhQvZni9GT3NVoknmoJCqeYJmA+CiDX
wZaBJHCJUh96qt7pZ1gYGnNycpXAbok2FCPKMdsIwZUw0c3+xc8DHK8rkr68QFMK
EjVpkVvQODacqy02ERpkCMKbHbg+uMkS/CMFPggwtWZ49oW3dpYkwKOMmvl5sx+l
pN+XsQ51xqKJEdP5tiUYhK+CaOPpXEXl/iJ2NVfzNNuoRzw8Q+NbDpvvXSkFtcln
oTr75/a8/XhZuHnEM83Pkq1yVJhzpDAf+GPeQk3uuo1gaF5Rl2pUsCwdMY5R80Cr
4UaJvT9Zu7H5f3abaQ1vLqV8KnFB4o/42+vLlRrvbBI3wmaXQ6py/WJxFwpTRa50
Xg+puvZvJSi0I3UNyyDvxtz0oM3bUfs976PtjQp6I/1no4Hy7lpnmc4390rLghWb
Dp+oUEliRAArufVUy9+hOP9k/UweaURYQxqOITtb3GmEl8IdRWJYmrIBqPJSxb7M
SOV6mC6V2FRU0/NDCLn+FxgMEq0cSBcjPswLB3jdFrt6xN8dRQGACAICljZpU8XJ
4Rda8Asr/KcBVquWwCnT8OPVCcOika1pw+QVRsY5zjySv5HA0oU9e/q2NoLXopED
tMUdwdK55ktbctt4Y/1MStpSVMbjbjbOHi+Q+ZYmvHFtAgNNIcE3/zJDgPXV1HfH
uYdfONKxVMi5ZQEODoLel6kanbJgcKmgQ1Sp5OfBC7PD32fTxdxrB7lPpThY2HVy
zwhnFe0PvljDxbrQMBSjasLvrmfBLjN/idL3RDQqAlP70CNFZ+OZXCs7L2DE9hOK
bofiH+GVXLg9cm5CjThIpGc3VuBnJ5ztp0RHmfomyvTVsZQ9tB5SqH/54BOAUcux
n83pVdmxsvykKk8Owu45OlbFnu4KoduLFr0jXO6ClI3ejmOQcUypuisAykwlE85Q
5yZrTvoMNn2JcR4yDPktTCPptFXo0I0rZWkRxe6LTUK1RAePBjYKxr9POoZx3mWf
khXGBaETeqmStJbDRJom7ocFl/dLCqzGKhBCGxNZgPJu1KIny78+6xiUr6fJTddZ
j0gu3oErhWfi1fCr8Ry8ZoEHljAVPaqmFjsg3MmbnEkW6tdm42As3C/W+WFzeGfH
ytUtJHM84KO+CkC4pN7ulAqhIgeBlC3yUNn2ZJ+hpycHgyYHCTrppRFuabUFMco1
ENF+3O8p1s05JILr9YSifpCCfiwS8KPpEw2LFcmMq5NHW5HJE88owh3WhYmrMM/7
3NKvF3LH8O/SCPlTr94JTeHYp6NtNpyYob8FrQ58rZJnw/9lbEnZ/YlgjeX+De1b
hhaZSyHrn7pddHiO8dG6KIuP/MLl5swswTrRtVSINjzkGqrMqyliWxwBGkXkaV9n
s/IAw1lzNkqsWB9i+wPN11lYxcZaXGvGMgdQRR4sxMUTptqQ3mzSxE7Jkm8JuzQy
QklR8iOrmeR9rv/cTaa0NaNSNSJN4Vrey9w7Pxqbec/lObuxwUaZvbENe1tlN9aO
PtuXwc0VvBKx6JN93qceqv9LpHk2mEoYr7iMZSGc0DsF4lM216eymN2zAxHL36vI
3tqRC5s8Yc62BOnJWGHuUXa9fdZaSbYe8Pl227Si34hCfwSAHlBZmdoCKtbEWQzw
Jia0bqS0wDS7CPgu4O+oUVFJSkS7lDn04aIc6lQERj2dEFOJJ+nJzrEwG4ePuOH4
PJ51IgQFB8P1ahFFTyJP1/HSDceL7ZhsT1tqjL6Tq8j8yUh66xdt2r7fhbQVqnQ/
qm5rgqN5hCZhONWjU9MGWH5RdioHgsSUGf+m4m8gYJuB+HpoGgFxtqZLketamoBB
1yB5n2VexnTNoBL9g6nIXNiaDl4ymZuuW5Zr+BEnN78eY4i5koGUVmmZbl2AgNIY
Zgov1Pp3FcQCcWoc07hPLpNDL2AdKPlerpNr60mr4PdmmwpdUvRMgFaLO9C9utns
17Xq0KW2gIWQhcuGT1BxP+oJh0AOudNYmrb2n2py5F064szmWj5S5Gh+Jf54yA3O
KbU/OSt4/B1Wck0sCJAAbEWthVT1Su7gqsB4+bRtHOriIjx0Q3CYKX4vCxO5RTHM
CrE8C0/Jw6z1+UQ6v9r3UU7WSXMjn2lkQzgg41nuzc/Nmj5s2/IYvWOK5vv0zQcj
buAamdIR4Cux6cWe98c7FwJDXAdlmQA1QpR0IPGohHi6RibACtEVcZFuhfiNuMju
53bMrJvacDVRBNUjwAsgJ09icm2IFnLixQxR/ImqKLFgiu7/Lm/t51pjhk1UJ9Th
1rriI5s/g0l10ZllqTYfLRJk81Q7F0LLSZza2lJnn+NM4I54J9We6Tdahzdq+WKe
sLwxSpgRlO65JsNSjMkoXyyHU2ISYBVXka1B6OdwOgWMoFrmk/6iL/Qjnbw2FbyP
SmqzcXOnTkt9P79ZSQuaN/XSSIS8MyDMsfIShqy1NKJmlDgNTrMx5W7tTQwkPjzI
5J8XKRpjfO37aa1/lXfBitmrMQNpgExQLmj1G50o4PeTIpuoGPNOk1Eov6KkzrrN
qn8g1c5YcMW40LCejbYrYHnzLIo9iSiuC3kjNFbggXEleTKQH0kfsodZ0GcFAxyp
SnnjAj5KCRJHJCJnv1vg+ZysbIanjgMV6tVhaymUBF9lQIBDQ/ZrdeOKHytNvdLL
gwRbHQuf9WHZfQpoh9QQ8+ZxXc0SnYq+cilB9Y3TbnyUqrM7/NZ6smT1hkyx03VF
W34y8HmtPuaUvgW/lw3tQFGPsg59qPfGd9xEQYqv0ADXBTxbsTV1s0F/+DGxSJYE
JewneqHdpv4x7bSZVfFSwoexAFcPmM6SlRaF+Jj2A0QoqfYFHawkiFq9Y68T5TV+
/17v5kNrnDviMAp8YwRouCDVRVow4QoIMoticJK3UEafbe5BYD6SZY7oXO5U8IN8
0KJOioAG7E+rHZey0uygXwzYZYjBjiX0LcbEoar2/Vdi4qqgazaCDV5u1MmhDiIH
5dvzjFd+/B6uST541ePOcINXrXuZ4CH5xsbbIIsSv0u9zeVOhj83xTUGhyYLJKj0
t0XF0fa7saQEo+88exYDEAK5Jog34tB7sj28i4k2mRz0IoVgqtTlVsp0sR+k2LH1
1/loIN4RXDkZpqqzL1d42zD+IpJ339W4CB8hAvlYYo7FyXDsbHTuhVaunGHiZaB7
igKqHgPtHWaaKwB+Nsl/OaF9jvczVtqDFCr+2jSFglDIXN0/3YVqULasvcyEHEVp
vBH37BZigE9YpMQj1xQ6keidAazAJ12Vy7dGMLgzCR70ZLUYK+96Vz4535N9eifM
k7hFZVGDff3qELUP14ZEzLCjxwnzjZko5oZLTX/xbIoFKJ4XB+0OUzOqe3vBw0Bn
IMOZ70bTEBieprnjXoUd2bqQobotEsbGhY4qHsOAB68Ivef5cyn5TkcTxonx9d+l
Pc8aWNi9C6FoDW38eZd4Nb+UlHTitTMuL9JeOMkBg3jwG7s6w6hcv4enGIiAaMYT
wJRyvCxOD/Ehiikp/VkNsHdrjN35sqyjlP3R5uoYE3inQrxzVDr5Ao8uhwSUaSvR
MdydIwn6djsJNLe/5eCQywio+spUlY6mYBNhjHkO7oKJuv8bJ7LD3mHlUdaI8Hi1
Ntm3lljQbZaeBXYjBKwWTO5FbAXBL7MaBI/XugQlq8b2mQkJeHaPyVYQTCuZ7Ace
MkDMZiBrCjFYvHWKvRNL66sPxtBnsf1KSwu/y2VlUu5qk4+BMB4GNVfFFRrGvKKD
LKOKTXBUqUUgCEokGWoe2z1kA098xEjYadymxraDeHWXW/gsbJWaJOUF4Wrtorel
4/ZPWyv0TDB0+0bXepe/zWizaIofIXVQRbUfuCKY9n1p8GRqHVH1jDIbC+mJWxqu
5s5i7SNzKWndF2Rzw1axYnTwaSi+aamA0QDDmuQbvhDxlHcwsiXl+aB6tSlV8H0P
vBqMTDnsi2UTzVORuC4fo9dnh0unVCIiSqJzPWKkdZa/y+KoTVt2sisVHzC4EfwA
LOFOLa19BWGM139uPjJf/cPVXUytaFLYtg/D35e5Iv6IAuc/fGbukRALLBNNIyot
TWtsMrnEgYm2TQmwHD8V/W42jCnCv75QCe/4RPIzUx8hfkKj2pawoJJEv+Apx6Cn
ftiV1d2FC2jqoIsz/o1HBkjqz/krjhTiHuzRF9CdRnbf8hnpPRqRrqRMeEJmEjUl
FCitBC3uC360wx9GW9qodvE5dWLRkuEL33AVoJnhLl9Bj2AR7JbmFusp8QISAi4o
XNY+gd+H6mqL2glmZuyMqNTtnTyFVD32bSlTmNT6JdPq6f1ZKdiazP7Ho0wrsor6
wNY3olw6Chb+freJjPr81go9Oe9QH4uVMo6nJM9XIScNSA5TQg3dWUEQU1B1FXii
6tiMrt6mUr98hAw26SF4TeDRrFKKBJiobSJfvSZs++2iWgkrSfEIiQj2jCgtqlq1
1+OsIjIaWDP/0niGUiqB/RW4Od9At1jJ1vtjeJ5BAmu5iwgbdZ2HXnDZiWAVmLuI
R5RrKvBZQ0YeJGKTESB3mATEAWMnO6h/7oMcE4R/D3MmOWx/tYhO54G5YoyzVfqn
yzya9OIaIsVgE+rcWmT5RuAC254uW/id2/IuE+YVYF3b/IPJxePkgPLp5FO7hT1Q
PB81/BSG10eeiSDI8HaUZ3PgyDzz4r3yYmLzjyUmFlCgEbgDURB8j5xblnBuXQ0z
0+iNOsm6WA2uLXt9BkwKec+U4xLZKHTferPu8jfOdhYXLXYD37fU5PyW/MpJb9dX
63qo1t4lyCOFqhuAPo5EF/PU9vpSfqdLmbv2yQHwkv4OMQfuzhajKxZNNehizzT2
2sOZKlvGc3U8+lnvJDK2dW06O91KaBI6XDIVJK1uWgvIV7rtAOufbllxFos8rNzu
jxO04cBXCNDWGX1dGC7KtX+VP81oo7/WylDquzeejRsemsfhwEWltWCd20P+aALt
3d6l+n3OV78YWEbXZAxvFsNt2y0Vjtq7VNK3/QsnKcZllb3PLlxLgZeLvnhwe5Iy
/U1P07t60nEbf2g/UeMWbzgkvwoPqix4r1SBGCg5MUh8L/bJK3lO7q7YM+vRzjsu
HUW9z5lhDTIOFqFZPaX0HPtwI355wmA37crFTv+h26bLKvaW5aZGPvp2HCMD3odL
Rot0L/NI4F34kbFhE6MxSW8to7Z7PQJPCZ1n92Jyk2kRftll3726rbOWsVYV7O6G
oQqghhx1eEyYvm7echHKknhBP7hQ3ujZ1zIp2p9jJjd4LKMSmdfMacC3ONfcd7XM
K8/ftz16xzyqGJUDOuGwfhss0KZx3M6OqU3QgR1cHAvHJXNFyMj97tVCZk7C1my7
40XYdpJ/YSt/031HUw0VfIS9+ydB0pdo7+TG98ZHMcX3/mEPBTrbgU2o8Wu9Mr4B
z59/PC1A1iqYFJ8v7H2KcBeD+C+IGKoWqG9/wu2U8F/bTTD0ORs71RK2lBrtiryn
JEApgDrOiwnBclhrHAr+3VLnzfEO+b21q/h+KkG0QTdQFMUcDRQEFW/7YxJj+xr2
n6j/G5avACBuDBUHrIfI3Q367XVlOv1qyX/7rQ45LceHtD5hDesEqmkYiF6seINr
0kGRDdlQw2VV9uBs5gTptLiZPv2t+9ak8/iM+Jt3XLYfz1PecK1C28saBacIcdOp
ytRnZw5AlFMgc1Xe9bB5N7SAnbmx6D3XYYca7Z9r0XeTZMT3X6BgarhvkCTCD7KB
I+/c2mNIbW9F93VTk8noMkSeq9zBc05i8QQRQ351hmpipN36jHxzUp/zu25Ns5X1
nz5ZVfnyARXsEtQA9RTFNMQKlbhljIYB0hLsa68F1QvtBWPUkuDtghpWtmI4ujBx
scSHJERZOrw3xZr2WiiM0ciy9ho+SwbzrCZ3v6Tlb6D9tu6PCpYwOiV8g/VaRMuP
r4mknw8mduwjEPI3ViVjAy/zxHSRB7TstL4Hy26E/6skRyAyJiws2cDOE8pHN+U2
yTo5LmjSOJbnM78xLSpiT2wn0K8bPQ+ii7MQ0dCfeYbGadW7071x5DhrGlcOdzvC
Kf758Dr7v9Uvyp71OO4RSqaWJF9mzO5RK197sy3fJSW+FfLdu9430+ckdX6i2zHD
6rLe3Ftyv/mXNyWqba5Oudl1gO44KCUqfB6zhb/bCE+VNvgXOsThXpP2tqqcVCQB
+824cs2HCsd14TfTRSalqLupQ0v3yPAZJ5Py8/BwcGRDWy8/KjMjpVWktB+jdCAf
c7CoM/TxYORpZvIBb47BLigtKk8fuXm+614Z1WZdpTFeRp6ISpMojLRjLIYFtSJN
pHK3d4JJKkoRHOiVJVvFgOD/g1H/eil8aiPPYxMvI9F9Ihakk/NZvrszgIWcTSdM
qeilb7Lap5Yvt114zIXNlgv+YyKI8jwQPi28Xh4fnnE1LxIAMm333jRjQ76lGoUp
PirOcVoe5FZJM7X0kY8gRCK0oK+ElQwF2isbpGIha8k8hvIRmGBUfi+vDn95S5Fh
rqqiygq1Tsv9OjISCvA481ovkUfwz+W3IBV8L5ku1NmDqrokL9qxDzFor50uEsdM
8Q3a9NSryHNPSheiLsUT2SILE3UZIqTwTpYmRa6wtPHxDn3akKeiIaoX0IVd6o5I
FRnwihVajWW+9XQ7B1bD51onKl9qIg/W0PEfWAT1WaoQRNMsMPHchd1ZgyZ48tuO
m5jH9JUJqYhlczUfPjV+adgUHttMbAhTNf72nlHMNGuh9ziNM3r1CBuuMj4pCyqG
`pragma protect end_protected
